magic
tech scmos
timestamp 1731366734
<< nwell >>
rect 0 50 204 88
rect 0 28 91 50
rect 167 49 204 50
<< ntransistor >>
rect 11 9 13 19
rect 56 9 58 19
rect 102 14 104 34
rect 119 14 121 34
rect 141 14 143 34
rect 158 14 160 34
rect 175 31 177 35
rect 191 31 193 35
<< ptransistor >>
rect 11 35 13 75
rect 33 35 35 75
rect 56 35 58 75
rect 78 35 80 75
rect 111 58 113 78
rect 150 58 152 78
rect 175 56 177 76
rect 191 56 193 76
<< ndiffusion >>
rect 10 9 11 19
rect 13 9 14 19
rect 55 9 56 19
rect 58 9 59 19
rect 101 14 102 34
rect 104 14 105 34
rect 118 14 119 34
rect 121 14 122 34
rect 140 14 141 34
rect 143 14 144 34
rect 157 14 158 34
rect 160 14 161 34
rect 174 31 175 35
rect 177 31 178 35
rect 190 31 191 35
rect 193 31 194 35
<< pdiffusion >>
rect 10 35 11 75
rect 13 35 14 75
rect 32 35 33 75
rect 35 35 36 75
rect 55 35 56 75
rect 58 35 59 75
rect 77 35 78 75
rect 80 35 81 75
rect 110 58 111 78
rect 113 58 114 78
rect 149 58 150 78
rect 152 58 153 78
rect 174 56 175 76
rect 177 56 178 76
rect 190 56 191 76
rect 193 56 194 76
<< ndcontact >>
rect 6 9 10 19
rect 14 9 19 19
rect 51 9 55 19
rect 59 9 64 19
rect 97 14 101 34
rect 105 14 110 34
rect 114 14 118 34
rect 122 14 127 34
rect 136 14 140 34
rect 144 14 149 34
rect 153 14 157 34
rect 161 14 166 34
rect 170 31 174 35
rect 178 31 182 35
rect 186 31 190 35
rect 194 31 198 35
<< pdcontact >>
rect 6 35 10 75
rect 14 35 18 75
rect 28 35 32 75
rect 36 35 40 75
rect 51 35 55 75
rect 59 35 63 75
rect 73 35 77 75
rect 81 35 85 75
rect 105 58 110 78
rect 114 58 118 78
rect 144 58 149 78
rect 153 58 157 78
rect 170 56 174 76
rect 178 56 182 76
rect 186 56 190 76
rect 194 56 198 76
<< polysilicon >>
rect 111 78 113 81
rect 150 78 152 81
rect 11 75 13 78
rect 33 75 35 78
rect 56 75 58 78
rect 78 75 80 78
rect 175 76 177 79
rect 191 76 193 79
rect 111 56 113 58
rect 150 56 152 58
rect 111 54 121 56
rect 150 54 160 56
rect 11 19 13 35
rect 33 14 35 35
rect 56 19 58 35
rect 78 14 80 35
rect 102 34 104 43
rect 119 42 121 54
rect 119 34 121 37
rect 141 34 143 43
rect 158 42 160 54
rect 158 34 160 37
rect 175 35 177 56
rect 191 35 193 56
rect 175 28 177 31
rect 191 28 193 31
rect 102 11 104 14
rect 119 10 121 14
rect 141 11 143 14
rect 158 10 160 14
rect 11 6 13 9
rect 56 6 58 9
<< polycontact >>
rect 97 37 102 42
rect 7 22 11 26
rect 29 14 33 19
rect 52 22 56 26
rect 74 14 78 19
rect 119 37 123 42
rect 137 37 141 42
rect 171 44 175 48
rect 158 37 162 42
rect 187 44 191 48
<< metal1 >>
rect 0 84 204 88
rect 6 75 10 84
rect 51 75 55 84
rect 114 78 119 84
rect 153 78 158 84
rect 18 35 19 75
rect 27 35 28 75
rect 14 30 32 35
rect 63 35 64 75
rect 72 35 73 75
rect 36 26 40 35
rect 59 30 77 35
rect 118 58 119 78
rect 157 58 158 78
rect 170 76 174 84
rect 186 76 190 84
rect 105 49 110 58
rect 105 45 123 49
rect 144 48 149 58
rect 178 48 182 56
rect 194 48 198 56
rect 144 45 171 48
rect 81 28 85 35
rect 105 34 110 45
rect 144 34 149 45
rect 178 45 187 48
rect 178 35 182 45
rect 194 44 204 48
rect 194 35 198 44
rect 0 22 7 26
rect 36 22 52 26
rect 6 5 10 9
rect 36 11 40 22
rect 19 9 40 11
rect 14 8 40 9
rect 51 5 55 9
rect 81 11 85 23
rect 64 9 85 11
rect 59 8 85 9
rect 97 11 101 14
rect 114 11 118 14
rect 97 8 118 11
rect 122 5 127 14
rect 136 11 140 14
rect 153 11 157 14
rect 136 8 157 11
rect 161 5 166 14
rect 170 5 174 31
rect 186 5 190 31
rect 0 0 204 5
<< m2contact >>
rect 69 14 74 19
<< metal2 >>
rect 128 46 158 49
rect 153 42 158 46
rect 114 28 119 37
rect 86 23 119 28
<< m123contact >>
rect 123 45 128 50
rect 92 37 97 42
rect 114 37 119 42
rect 132 37 137 42
rect 153 37 158 42
rect 81 23 86 28
rect 24 14 29 19
<< metal3 >>
rect 92 57 135 61
rect 92 42 97 57
rect 132 42 135 57
rect 92 19 96 37
rect 0 14 24 19
rect 29 14 96 19
<< labels >>
rlabel metal1 2 23 2 23 3 d
rlabel metal3 1 16 1 16 3 Clk
rlabel metal2 88 25 88 25 1 qq
rlabel metal1 79 2 79 2 1 gnd
rlabel metal1 76 85 76 85 5 vdd
rlabel metal1 45 24 45 24 1 l1
rlabel metal1 163 46 163 46 1 q_preinv
rlabel metal1 201 46 201 46 7 q
<< end >>
