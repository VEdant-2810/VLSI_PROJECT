
.include all_subckts.spice

Vdd vdd gnd {SUPPLY}

Vclk clk 0 PULSE(0 {SUPPLY} 2n 100p 100p 30n 60n)
Vd   D   0 PULSE(0 {SUPPLY} 1n 100p 100p 9n 18n)  
*D is delayed by 5ns, for setup time and holdtime violation protection  


Xff1 clk D Q vdd gnd ff_1bit 

Cq Q gnd 10f

.tran 1n 340n 

.control
run

meas tran Q_delay_fall TRIG v(clk) VAL=0.9 RISE=3 TARG v(Q) val=0.9 FALL=1
meas tran Q_delay_rise TRIG v(clk) VAL=0.9 RISE=4 TARG v(Q) VAL=0.9 RISE=1
let tp2q = (Q_delay_rise + Q_delay_fall)/2
print tp2q;

meas tran tsu_r TRIG v(D) VAL=0.9 RISE=4 TARG v(Xff1.A) VAL=0.9 FALL=3
meas tran tsu_f TRIG v(D) VAL=0.9 FALL=3 TARG v(Xff1.A) VAL=0.9 RISE=2
let tsu = (tsu_r + tsu_f)/2
print tsu;


plot V(D)+4 V(clk)+2 V(Q) V(Xff1.A)+6
.endc
.end