magic
tech scmos
timestamp 1764705872
use nmos  nmos_2 ~/Documents/magiccccccc
timestamp 1764668464
transform -1 0 66 0 1 -4
box -10 -25 20 -5
use nmos  nmos_1
timestamp 1764668464
transform 1 0 9 0 1 -44
box -10 -25 20 -5
use nmos  nmos_0
timestamp 1764668464
transform 1 0 10 0 1 -16
box -10 -25 20 -5
use pmos  pmos_0 ~/Documents/magiccccccc
timestamp 1764668421
transform 1 0 10 0 1 11
box -10 -11 20 18
<< labels >>
rlabel space 2 -24 2 -24 3 gi
rlabel space 72 -27 72 -27 7 ci
rlabel space 74 -13 74 -13 7 pi
rlabel metal1 -13 -25 -13 -25 3 clk
rlabel metal1 28 -12 28 -12 1 out
rlabel space 12 26 12 26 5 vdd!
rlabel space 13 -67 13 -67 1 gnd!
<< end >>
