magic
tech scmos
timestamp 1764806298
<< nwell >>
rect 462 353 463 356
rect 928 355 929 356
<< metal1 >>
rect 1182 364 1248 365
rect 1182 363 1252 364
rect 1164 362 1252 363
rect -6 358 44 360
rect 1164 358 1186 362
rect -6 355 50 358
rect 0 353 50 355
rect 174 354 380 357
rect 463 356 668 357
rect 1095 356 1176 358
rect 462 354 668 356
rect 462 353 463 354
rect 564 352 667 354
rect 758 353 964 356
rect 1062 355 1176 356
rect 1053 352 1176 355
rect 1373 361 1472 366
rect 85 265 91 285
rect 375 255 379 286
rect 668 245 675 283
rect 966 248 971 283
rect 1286 252 1291 293
rect 1463 212 1472 361
rect -34 195 77 200
rect -120 163 -103 167
rect -159 139 -145 143
rect -141 -32 -134 125
rect -34 10 -27 195
rect 890 193 958 198
rect 1272 175 1294 180
rect 1315 175 1374 179
rect -3 122 5 169
rect 40 170 45 174
rect 112 170 383 171
rect 40 167 98 170
rect 112 168 388 170
rect 402 168 433 171
rect 1272 170 1277 175
rect 117 167 388 168
rect 40 123 45 167
rect 428 152 433 168
rect 656 166 679 170
rect 699 166 973 170
rect 993 166 1277 170
rect 656 152 662 166
rect 428 150 662 152
rect 1276 152 1292 155
rect 428 148 660 150
rect 86 143 90 147
rect 373 146 377 147
rect 369 143 377 146
rect 671 145 672 146
rect 369 134 373 143
rect 658 142 672 145
rect 954 142 968 146
rect 658 141 673 142
rect 283 129 373 134
rect 658 135 662 141
rect 590 131 662 135
rect 954 133 958 142
rect 1276 141 1280 152
rect 1184 136 1281 141
rect 1368 139 1374 175
rect 1464 143 1471 212
rect 1399 139 1472 143
rect 883 128 958 133
rect -4 119 6 122
rect 30 118 45 123
rect 150 108 157 121
rect 47 104 50 107
rect 46 98 50 104
rect 150 104 329 108
rect 441 107 447 124
rect 734 122 741 123
rect 731 108 741 122
rect 1032 116 1039 123
rect 1349 119 1355 131
rect 1032 109 1241 116
rect 1349 115 1375 119
rect 1402 115 1451 119
rect 150 103 185 104
rect -14 94 5 98
rect 33 94 50 98
rect -14 91 1 94
rect 441 102 630 107
rect 731 103 922 108
rect 1032 106 1039 109
rect -14 10 -7 91
rect 17 20 24 80
rect 67 64 86 67
rect 372 64 378 68
rect 56 36 87 40
rect 1201 43 1287 48
rect 303 36 374 40
rect 46 10 51 24
rect 61 22 66 36
rect 657 35 667 39
rect 925 35 963 39
rect 657 30 663 35
rect 610 23 662 30
rect 1244 12 1286 16
rect -34 8 91 10
rect -34 6 87 8
rect -34 0 -27 6
rect -86 -32 -32 -27
rect -160 -38 -32 -32
rect -160 -224 -155 -38
rect -86 -39 -32 -38
rect -14 -125 -7 6
rect 329 5 373 9
rect 629 4 669 8
rect 902 4 969 8
rect 1372 2 1376 104
rect 1253 -3 1289 2
rect 1309 -2 1377 2
rect 29 -11 89 -6
rect 108 -10 378 -6
rect 399 -10 669 -6
rect 694 -13 964 -6
rect 1253 -7 1258 -3
rect 988 -11 1258 -7
rect 1072 -66 1097 -62
rect 1125 -66 1202 -62
rect 1157 -67 1202 -66
rect 778 -76 808 -72
rect 836 -76 912 -71
rect 156 -92 185 -88
rect 213 -91 285 -88
rect 489 -89 514 -85
rect 543 -89 620 -86
rect 574 -90 620 -89
rect -14 -145 -8 -125
rect 278 -157 285 -91
rect 613 -158 620 -90
rect 900 -148 911 -76
rect 1197 -135 1202 -67
rect 871 -170 883 -169
rect -96 -175 -59 -172
rect 67 -176 251 -172
rect 240 -180 251 -176
rect 559 -173 564 -172
rect 559 -177 588 -173
rect 709 -176 883 -170
rect 709 -177 871 -176
rect 559 -178 564 -177
rect 366 -182 564 -178
rect 995 -180 1177 -176
rect -18 -204 -10 -188
rect -162 -239 -155 -224
rect -23 -206 -10 -204
rect -162 -299 -156 -239
rect -23 -243 -15 -206
rect 65 -248 131 -244
rect 272 -249 281 -198
rect 616 -245 620 -191
rect 709 -247 750 -243
rect 904 -246 910 -195
rect 366 -254 418 -249
rect 995 -250 1036 -246
rect 1197 -250 1202 -198
rect 1292 -254 1313 -250
rect -162 -313 -155 -299
<< m2contact >>
rect -6 345 0 355
rect 281 348 287 354
rect 575 346 581 352
rect 870 345 876 353
rect 1192 351 1198 362
rect -7 255 -1 261
rect 85 259 91 265
rect 281 255 286 260
rect 375 247 382 255
rect 575 254 581 260
rect 870 253 876 259
rect 668 237 675 245
rect 1192 263 1197 270
rect 966 239 971 248
rect 1286 242 1291 252
rect 1190 221 1197 228
rect 1366 220 1374 226
rect 169 211 176 218
rect 279 213 286 220
rect 455 211 463 218
rect 581 208 589 215
rect 749 210 757 217
rect 876 208 884 215
rect 1044 210 1051 217
rect 77 195 85 200
rect -103 163 -92 170
rect -117 136 -109 145
rect 958 193 967 199
rect 890 185 900 193
rect -4 169 5 178
rect 88 137 95 143
rect 275 129 283 136
rect 378 138 385 143
rect 582 130 590 137
rect 673 136 678 142
rect 968 136 973 142
rect 1289 144 1295 151
rect 874 128 883 133
rect 1179 128 1191 136
rect -14 98 -6 104
rect 157 92 168 103
rect 489 89 498 102
rect 778 90 787 103
rect 1072 97 1083 109
rect 1284 76 1290 83
rect 86 68 92 73
rect 374 68 381 73
rect 669 67 674 73
rect 964 67 969 73
rect 1201 48 1210 57
rect 48 36 56 41
rect 296 36 303 45
rect 17 13 24 20
rect 918 35 925 41
rect 602 23 610 31
rect 1231 12 1244 19
rect -32 -35 -23 -25
rect 321 5 329 10
rect 618 4 629 10
rect 891 4 902 9
rect 1399 100 1414 108
rect 24 -13 29 -3
rect 1072 -62 1081 -53
rect 778 -72 787 -63
rect 156 -88 165 -81
rect 489 -85 498 -78
rect -16 -157 -7 -145
rect 278 -166 286 -157
rect 613 -164 620 -158
rect 904 -162 912 -148
rect 1197 -156 1202 -135
rect -107 -179 -96 -172
rect -17 -188 -9 -180
rect 278 -198 286 -189
rect 614 -191 620 -183
rect 906 -195 912 -185
rect 1197 -198 1202 -188
rect -85 -273 -79 -267
rect -155 -322 -148 -305
rect -109 -319 -104 -313
rect 54 -320 64 -311
rect 189 -324 194 -319
rect 362 -322 367 -317
rect 534 -319 539 -314
rect 707 -317 712 -312
rect 820 -322 825 -317
rect 992 -320 997 -315
rect 1114 -326 1119 -321
<< metal2 >>
rect -6 261 0 345
rect -67 172 -4 176
rect -68 169 -4 172
rect -68 168 -57 169
rect -92 163 -57 168
rect -109 136 -95 143
rect -68 50 -57 163
rect 36 159 41 231
rect 85 196 91 259
rect 281 260 286 348
rect 575 260 581 346
rect 870 259 875 345
rect 1192 270 1198 351
rect 176 213 279 218
rect 323 211 328 231
rect 296 207 328 211
rect -45 155 41 159
rect -68 49 -56 50
rect -67 -71 -56 49
rect -45 41 -39 155
rect 88 136 95 137
rect 73 132 275 136
rect 88 129 275 132
rect -14 104 -6 110
rect 51 49 56 118
rect 88 73 93 129
rect 51 45 77 49
rect -45 36 48 41
rect 18 -25 24 13
rect -23 -35 24 -25
rect 18 -36 24 -35
rect -120 -73 -56 -71
rect -120 -78 -57 -73
rect -115 -179 -107 -78
rect 73 -115 77 45
rect 156 -81 167 92
rect 296 45 300 207
rect 374 200 381 247
rect 1285 242 1286 243
rect 618 224 622 230
rect 602 223 622 224
rect 602 221 621 223
rect 463 211 581 214
rect 315 195 381 200
rect 315 5 321 195
rect 378 134 382 138
rect 378 130 582 134
rect 339 -58 343 118
rect 378 73 382 130
rect 338 -78 343 -58
rect 334 -85 343 -78
rect 489 -78 498 89
rect 602 31 606 221
rect 669 200 675 237
rect 757 210 876 213
rect 614 193 675 200
rect 614 4 618 193
rect 671 132 676 136
rect 671 128 874 132
rect 635 45 639 117
rect 671 73 676 128
rect 635 -6 640 45
rect 636 -78 640 -6
rect 778 -63 788 90
rect 891 9 897 185
rect 913 35 918 230
rect 967 194 971 239
rect 1167 226 1173 227
rect 1167 221 1190 226
rect 1235 221 1239 239
rect 1167 215 1173 221
rect 1051 210 1173 215
rect 1201 217 1239 221
rect 1201 201 1206 217
rect 1285 208 1291 242
rect 1374 220 1450 226
rect 1280 207 1291 208
rect 1238 206 1294 207
rect 1224 203 1294 206
rect 966 132 972 136
rect 966 128 1179 132
rect 930 48 934 117
rect 966 73 972 128
rect 930 -6 935 48
rect 334 -106 342 -85
rect 636 -90 639 -78
rect 931 -87 935 -6
rect 1072 -53 1083 97
rect 1201 57 1207 201
rect 1224 138 1234 203
rect 1238 202 1294 203
rect 1272 201 1294 202
rect 1224 8 1231 138
rect 1250 -56 1254 126
rect 1286 83 1292 144
rect 1438 105 1448 220
rect 1414 99 1448 105
rect 1438 98 1448 99
rect 1205 -67 1255 -56
rect 636 -96 654 -90
rect -74 -123 77 -115
rect 335 -117 342 -106
rect 643 -103 654 -96
rect 856 -91 935 -87
rect 1151 -87 1154 -85
rect 1213 -87 1224 -67
rect 856 -94 1023 -91
rect 1151 -94 1225 -87
rect 856 -96 934 -94
rect 643 -109 655 -103
rect -101 -186 -97 -179
rect -101 -189 -79 -186
rect -82 -267 -79 -189
rect -73 -202 -65 -123
rect 73 -124 77 -123
rect 226 -123 342 -117
rect 570 -113 657 -109
rect -17 -180 -10 -157
rect 226 -208 230 -123
rect 279 -189 285 -166
rect 570 -203 574 -113
rect 614 -183 620 -164
rect 856 -210 859 -96
rect 906 -185 912 -162
rect 1151 -210 1154 -94
rect 1182 -95 1220 -94
rect 1197 -188 1202 -156
rect -148 -318 -109 -314
rect 64 -319 147 -315
rect 64 -320 189 -319
rect 106 -324 189 -320
rect 712 -317 773 -313
rect 759 -318 773 -317
rect 367 -323 537 -319
rect 759 -322 820 -318
rect 997 -320 1110 -317
rect 1107 -323 1110 -320
rect 1107 -326 1114 -323
<< m3contact >>
rect -95 134 -85 145
rect 73 136 81 143
rect -14 110 -6 118
<< metal3 >>
rect -85 136 73 142
rect -81 110 -14 118
use 1bit_mcl  1bit_mcl_0
timestamp 1764797379
transform 1 0 57 0 1 104
box -71 -114 174 253
use inverter  inverter_0
timestamp 1764702656
transform 1 0 13 0 1 104
box -10 -25 20 18
use xorg  xorg_0
timestamp 1764782750
transform 1 0 -61 0 1 -201
box -62 -125 143 29
use 1bit_mcl  1bit_mcl_1
timestamp 1764797379
transform 1 0 344 0 1 104
box -71 -114 174 253
use inverter  inverter_2
timestamp 1764702656
transform 1 0 193 0 1 -82
box -10 -25 20 18
use xorg  xorg_1
timestamp 1764782750
transform 1 0 238 0 1 -207
box -62 -125 143 29
use 1bit_mcl  1bit_mcl_2
timestamp 1764797379
transform 1 0 639 0 1 103
box -71 -114 174 253
use inverter  inverter_3
timestamp 1764702656
transform 1 0 524 0 1 -79
box -10 -25 20 18
use xorg  xorg_2
timestamp 1764782750
transform 1 0 582 0 1 -202
box -62 -125 143 29
use inverter  inverter_4
timestamp 1764702656
transform 1 0 816 0 1 -66
box -10 -25 20 18
use xorg  xorg_3
timestamp 1764782750
transform 1 0 868 0 1 -205
box -62 -125 143 29
use 1bit_mcl  1bit_mcl_3
timestamp 1764797379
transform 1 0 934 0 1 103
box -71 -114 174 253
use inverter  inverter_5
timestamp 1764702656
transform 1 0 1105 0 1 -56
box -10 -25 20 18
use xorg  xorg_4
timestamp 1764782750
transform 1 0 1163 0 1 -209
box -62 -125 143 29
use 1bit_mcl  1bit_mcl_4
timestamp 1764797379
transform 1 0 1255 0 1 112
box -71 -114 174 253
use inverter  inverter_1
timestamp 1764702656
transform 1 0 1382 0 1 125
box -10 -25 20 18
use inverter  inverter_6
timestamp 1764702656
transform 1 0 -137 0 1 149
box -10 -25 20 18
<< labels >>
rlabel metal1 157 167 165 169 1 vff
rlabel metal1 157 167 165 169 1 vdd
rlabel metal1 161 -9 169 -7 1 gnd
rlabel space 1289 151 1293 154 1 clk
rlabel space 85 37 88 39 1 A0
rlabel space 87 6 90 8 1 B0
rlabel space 50 229 53 231 1 A0
rlabel space 70 289 76 292 1 B0
rlabel metal1 198 105 204 108 1 C0bar
rlabel space 374 36 380 39 1 A1
rlabel space 374 6 380 9 1 B1
rlabel space 335 230 341 233 1 A1
rlabel space 357 289 363 292 1 B1
rlabel metal1 501 102 507 105 1 C1bar
rlabel space 668 36 674 39 1 A2
rlabel space 668 5 674 8 1 B2
rlabel space 632 229 638 232 1 A2
rlabel space 653 288 659 291 1 B2
rlabel metal1 823 104 829 107 1 C2bar
rlabel space 965 35 971 38 1 A3
rlabel space 964 4 970 7 1 B3
rlabel space 927 228 933 231 1 A3
rlabel space 948 289 954 292 1 B3
rlabel metal1 1105 111 1111 114 1 C3bar
rlabel space 1285 45 1291 48 1 A4
rlabel space 1285 13 1291 16 1 B4
rlabel space 1249 237 1255 240 1 A4
rlabel space 1279 291 1285 294 1 B4
rlabel space 1340 127 1346 130 1 Coutbar
rlabel metal1 1417 117 1427 118 1 Cout
rlabel metal2 73 -123 76 -105 1 P0
rlabel metal2 988 -94 1019 -91 1 P3
rlabel metal1 93 -248 110 -244 1 S0
rlabel metal1 391 -254 400 -251 1 S1
rlabel metal2 1218 -66 1233 -59 1 P4
rlabel metal1 726 -246 742 -244 1 S2
rlabel metal1 1015 -250 1031 -248 1 S3
rlabel metal1 1300 -254 1310 -252 1 S4
rlabel metal2 323 -121 334 -119 1 P1
rlabel metal2 646 -108 648 -101 1 P2
rlabel metal1 62 23 63 27 1 A0
rlabel metal1 48 14 49 18 1 B0
rlabel metal1 349 36 355 38 1 A1
rlabel metal1 350 5 356 7 1 B1
rlabel metal1 651 24 657 26 1 A2
rlabel metal1 646 6 652 8 1 B2
rlabel metal1 944 35 950 37 1 A3
rlabel metal1 940 5 946 7 1 B3
rlabel metal1 1264 44 1270 46 1 A4
rlabel metal1 1261 13 1267 15 1 B4
rlabel metal2 -105 137 -97 139 1 clk_mca
rlabel metal1 -156 139 -152 142 1 clk
rlabel metal3 -80 111 -76 114 1 Cin
<< end >>
