magic
tech scmos
timestamp 1731343607
<< nwell >>
rect -23 38 65 113
<< ntransistor >>
rect -12 19 -10 29
rect 9 19 11 29
rect 30 19 32 29
rect 52 19 54 29
<< ptransistor >>
rect -12 45 -10 105
rect 9 45 11 105
rect 30 45 32 105
rect 52 45 54 65
<< ndiffusion >>
rect -13 19 -12 29
rect -10 19 -9 29
rect 8 19 9 29
rect 11 19 12 29
rect 29 19 30 29
rect 32 19 33 29
rect 51 19 52 29
rect 54 19 55 29
<< pdiffusion >>
rect -13 45 -12 105
rect -10 45 -9 105
rect 8 45 9 105
rect 11 45 12 105
rect 29 45 30 105
rect 32 45 33 105
rect 51 45 52 65
rect 54 45 55 65
<< ndcontact >>
rect -18 19 -13 29
rect -9 19 -4 29
rect 3 19 8 29
rect 12 19 17 29
rect 25 19 29 29
rect 33 19 38 29
rect 47 19 51 29
rect 55 19 59 29
<< pdcontact >>
rect -17 45 -13 105
rect -9 45 -5 105
rect 4 45 8 105
rect 12 45 16 105
rect 25 45 29 105
rect 33 45 37 105
rect 47 45 51 65
rect 55 45 59 65
<< polysilicon >>
rect -12 105 -10 108
rect 9 105 11 108
rect 30 105 32 108
rect 52 65 54 68
rect -12 29 -10 45
rect 9 29 11 45
rect 30 29 32 45
rect 52 29 54 45
rect -12 16 -10 19
rect 9 16 11 19
rect 30 16 32 19
rect 52 16 54 19
<< polycontact >>
rect -16 32 -12 36
rect 5 32 9 36
rect 26 32 30 36
rect 47 32 52 37
<< metal1 >>
rect -23 109 65 113
rect -17 105 -13 109
rect -5 45 -4 105
rect 3 45 4 105
rect -9 40 8 45
rect 16 45 17 105
rect 24 45 25 105
rect 12 40 29 45
rect 47 65 51 109
rect -20 32 -16 36
rect 1 32 5 36
rect 22 32 26 36
rect 55 36 59 45
rect 55 32 65 36
rect 55 29 59 32
rect -18 15 -13 19
rect 3 15 8 19
rect 25 15 29 19
rect 47 15 51 19
rect -23 10 65 15
<< metal2 >>
rect 33 37 38 40
rect 33 34 42 37
rect -4 29 12 34
rect 17 29 33 34
rect 38 32 42 34
<< m123contact >>
rect 33 40 38 45
rect -9 29 -4 34
rect 12 29 17 34
rect 33 29 38 34
rect 42 32 47 37
<< labels >>
rlabel metal1 62 33 63 34 7 out
rlabel metal1 46 12 47 13 1 gnd
rlabel metal1 -19 33 -18 34 3 aa
rlabel metal1 24 35 24 35 1 cc
rlabel metal2 40 34 40 34 1 ee
rlabel metal1 32 111 33 112 5 vdd
rlabel metal1 3 35 3 35 1 bb
<< end >>
