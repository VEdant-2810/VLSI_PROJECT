* SPICE3 file created from manch.ext - technology: scmos
.include TSMC_180nm.txt
.option scale=0.09u

M1000 out G X Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1001 X clk gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1002 out P Cin Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1003 out clk vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=40 ps=26

C0 out clk 0.05fF
C1 X G 0.05fF
C2 P Cin 0.05fF
C3 X clk 0.05fF
C4 vdd vdd 0.08fF
C5 gnd X 0.08fF
C6 out P 0.05fF
C7 vdd clk 0.07fF
C8 out X 0.08fF
C9 vdd out 0.03fF
C10 out G 0.05fF
C11 out Cin 0.08fF
C12 out vdd 0.12fF
C13 gnd clk 0.05fF
C14 vdd Gnd 0.03fF
C15 vdd Gnd 0.58fF
C16 out Gnd 0.32fF
C17 Cin Gnd 0.11fF
C18 P Gnd 0.16fF
C19 X Gnd 0.22fF
C20 gnd Gnd 0.11fF
C21 clk Gnd 0.55fF
C22 G Gnd 0.16fF

Vclk clk 0 PULSE(0 1.8 0 100p 100p 5n 10n)
Vc Cin 0 PULSE(0 1.8 0 100p 100p 4n 8n)
Vdd vdd 0 1.8


