* SPICE3 file created from nandg.ext - technology: scmos

.option scale=0.09u

M1000 m1_30_1# A m1_26_n48# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 m1_26_n48# m1_54_n51# nmos_1/a_n1_n17# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1002 m1_30_1# A vdd pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=80 ps=52
M1003 m1_30_1# m1_54_n51# vdd pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
