

.include all_subckts.spice
Vdd vdd gnd {SUPPLY}

Vclk clk 0 PULSE(0 {SUPPLY} 10n 100p 100p 10n 20n)

Va A 0 PULSE(0 {SUPPLY} 80n 100p 100p 80n 160n)
Vb B 0 PULSE(0 {SUPPLY} 40n 100p 100p 40n 80n)
Vc Cin 0 PULSE(0 {SUPPLY} 20n 100p 100p 20n 40n)

C_cinbar Cinbar gnd 10f
Xcin_p Cinbar Cin vdd vdd pmos wp={1.8u}
Xcin_n Cinbar Cin gnd gnd nmos wn={0.9u}


Xmcl clk A B Cin Cinbar Cout Coutbar Sum vdd gnd mcl
C_cout Cout gnd 10f
C_coutbar Coutbar gnd 10f
C_sum Sum gnd 10f

.tran 1n 320n 

.control
run
plot V(A) V(B)+2 V(Cin)+4 V(Cout)+6 V(Sum)+8 V(clk)+10
.endc
.end
