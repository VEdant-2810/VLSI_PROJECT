.include 'TSMC_180nm.txt'

.option scale=0.09u
.global gnd vdd


M1000 a_362_217 clk a_355_217 0 CMOSN w=20 l=2 ad=100 pd=50 as=2550 ps=1290
M1001 a_362_217 a_310_170 vdd vdd CMOSP w=40 l=2 ad=200 pd=90 as=18800 ps=8930
M1002 X D vdd vdd CMOSP w=40 l=2 ad=400 pd=190 as=0 ps=0
M1003 a_310_170 a_258_170 0 0 CMOSN w=20 l=2 ad=100 pd=50 as=32400 ps=1800
M1004 a_407_217 a_362_217 0 0 CMOSN w=20 l=2 ad=200 pd=100 as=0 ps=0
M1005 a_459_241 a_414_217 0 0 CMOSN w=20 l=2 ad=100 pd=50 as=200 ps=100

M1006 Q a_459_241 vdd vdd CMOSP w=40 l=2 ad=200 pd=90 as=32400 ps=1620

M1007 a_310_170 clk a_303_211 vdd CMOSP w=40 l=2 ad=200 pd=90 as=32400 ps=1620
M1008 a_258_170 D 0 0 CMOSN w=20 l=2 ad=100 pd=50 as=0 ps=0
M1009 a_355_217 a_310_170 0 0 CMOSN w=20 l=2 ad=0 pd=0 as=0 ps=0
M1010 a_258_170 clk X vdd CMOSP w=40 l=2 ad=200 pd=90 as=0 ps=0
M1011 a_459_241 a_414_217 vdd vdd CMOSP w=40 l=2 ad=200 pd=90 as=0 ps=0

M1012 a_414_217 clk a_407_217 0 CMOSN w=20 l=2 ad=100 pd=50 as=0 ps=0
M1013 Q a_459_241 0 0 CMOSN w=20 l=2 ad=100 pd=50 as=0 ps=0

M1014 a_303_211 a_258_170 vdd vdd CMOSP w=40 l=2 ad=0 pd=0 as=0 ps=0
M1015 a_414_217 a_362_217 vdd vdd CMOSP w=40 l=2 ad=200 pd=90 as=0 ps=0

C0 a_459_241 0 0.32fF
C1 a_310_170 clk 0.11fF
C2 a_407_217 a_362_217 0.13fF
C3 a_414_217 a_362_217 0.08fF
C4 a_303_211 vdd 0.71fF
C5 D X 0.13fF
C6 X vdd 0.71fF
C7 D a_258_170 0.08fF
C8 0 a_362_217 0.06fF
C9 a_310_170 a_362_217 0.08fF
C10 a_362_217 clk 0.11fF
C11 vdd Q 0.58fF
C12 a_258_170 vdd 0.34fF
C13 a_414_217 vdd 0.60fF
C14 a_258_170 a_303_211 0.13fF
C15 a_459_241 Q 0.08fF
C16 0 D 0.06fF
C17 0 Q 0.26fF
C18 X a_258_170 0.50fF
C19 D clk 0.25fF
C20 a_310_170 vdd 0.30fF
C21 clk vdd 0.35fF
C22 a_407_217 a_414_217 0.23fF
C23 a_310_170 a_303_211 0.50fF
C24 a_303_211 clk 0.05fF
C25 0 a_355_217 0.23fF
C26 a_414_217 vdd 0.10fF
C27 a_310_170 a_355_217 0.13fF
C28 clk a_355_217 0.05fF
C29 X clk 0.05fF
C30 0 a_258_170 0.29fF
C31 a_407_217 0 0.23fF
C32 a_459_241 a_414_217 0.08fF
C33 a_310_170 a_258_170 0.08fF
C34 a_258_170 clk 0.36fF
C35 a_362_217 vdd 0.82fF
C36 a_407_217 clk 0.05fF
C37 0 a_414_217 0.06fF
C38 a_414_217 clk 0.08fF
C39 a_459_241 vdd 0.68fF
C40 a_362_217 a_355_217 0.23fF
C41 0 a_310_170 0.29fF
C42 0 clk 0.16fF
C43 D vdd 0.25fF
C44 0 0 0.51fF
C45 a_407_217 0 0.19fF
C46 a_355_217 0 0.19fF
C47 0 0 0.45fF
C48 clk 0 0.62fF
C49 Q 0 0.11fF
C50 a_303_211 0 0.00fF
C51 X 0 0.00fF
C52 a_362_217 0 0.79fF
C53 a_310_170 0 0.12fF
C54 a_258_170 0 0.52fF
C55 D 0 0.38fF
C56 a_459_241 0 0.32fF
C57 a_414_217 0 0.41fF
C58 vdd 0 2.48fF
C59 vdd 0 0.43fF
.ic v(a_414_217)=0 v(Q)=0

.tran 0.1ns 100ns

Vsupply vdd 0 1.8
Vclk clk 0 PULSE(0 1.8 1ns 100ps 100ps 10ns 20ns)
Vdata D 0 PULSE(0 1.8 0ns 100ps 100ps 4ns 8ns)

.control
    run

    meas tran tcq_rise TRIG v(clk) VAL=0.9 RISE=3 TARG v(Q) VAL=0.9 RISE=2
    meas tran tcq_fall TRIG v(clk) VAL=0.9 RISE=4 TARG v(Q) VAL=0.9 FALL=2

    let delay = (tcq_rise + tcq_fall)/2
    print delay


    meas tran tsu_rise TRIG v(D) VAL=0.9 FALL=3  TARG v(X) VAL=1.4 RISE=3
    meas tran tsu_fall TRIG v(D) VAL=0.9 RISE=3 TARG v(X) VAL=1.4 FALL=3

    let tsu = (tsu_rise+ tsu_fall)/2
    print tsu

    plot v(clk)+4 v(D)+2 v(Q)-2 v(X)
.endc
