magic
tech scmos
timestamp 1731573344
<< nwell >>
rect -290 169 -87 173
rect -63 169 137 173
rect -290 135 -86 169
rect -290 113 -199 135
rect -123 134 -86 135
rect -67 135 137 169
rect -67 113 24 135
rect 100 134 137 135
rect 388 130 592 168
rect 388 108 479 130
rect 555 129 592 130
rect 218 89 245 90
rect -290 41 -86 79
rect -290 19 -199 41
rect -123 40 -86 41
rect 2 28 26 63
rect 32 60 65 68
rect 188 65 245 89
rect 32 36 89 60
rect 212 57 245 65
rect 251 62 275 97
rect 320 89 347 90
rect 290 65 347 89
rect 314 57 347 65
rect 353 62 377 97
rect 32 35 59 36
rect 95 2 179 57
rect 398 34 602 72
rect 219 17 246 18
rect 109 0 121 2
rect 189 -7 246 17
rect -290 -53 -86 -15
rect -290 -75 -199 -53
rect -123 -54 -86 -53
rect 48 -73 83 -8
rect 213 -15 246 -7
rect 252 -10 276 25
rect 320 17 347 18
rect 290 -7 347 17
rect 314 -15 347 -7
rect 353 -10 377 25
rect 398 12 489 34
rect 565 33 602 34
rect -290 -146 -86 -108
rect -17 -113 7 -78
rect 13 -81 60 -73
rect 93 -79 161 -44
rect 179 -77 263 -22
rect 273 -77 357 -22
rect 367 -26 437 -22
rect 451 -26 655 -19
rect 367 -57 655 -26
rect 367 -77 542 -57
rect 618 -58 655 -57
rect 451 -79 542 -77
rect 13 -105 70 -81
rect 13 -106 40 -105
rect -290 -168 -199 -146
rect -123 -147 -86 -146
rect -290 -240 -86 -202
rect 29 -214 64 -149
rect 93 -166 190 -132
rect 204 -163 273 -128
rect 347 -211 402 -145
rect 437 -152 528 -130
rect 604 -152 641 -151
rect 437 -190 641 -152
rect -290 -262 -199 -240
rect -123 -241 -86 -240
rect -34 -254 -10 -219
rect -4 -220 64 -214
rect -4 -246 53 -220
rect -4 -247 23 -246
rect 101 -265 198 -231
rect 204 -247 292 -212
rect -290 -334 -86 -296
rect -290 -356 -199 -334
rect -123 -335 -86 -334
rect 12 -355 47 -290
rect -290 -428 -86 -390
rect -52 -395 -28 -360
rect -22 -363 25 -355
rect -22 -387 35 -363
rect 105 -366 193 -331
rect 204 -341 297 -306
rect 347 -310 422 -223
rect 440 -288 500 -197
rect 440 -331 478 -288
rect 349 -364 478 -331
rect -22 -388 5 -387
rect -290 -450 -199 -428
rect -123 -429 -86 -428
rect -6 -496 29 -431
rect 98 -460 163 -425
rect 204 -435 269 -400
rect 349 -401 479 -364
rect 349 -442 444 -401
<< ntransistor >>
rect -279 94 -277 104
rect -234 94 -232 104
rect -188 99 -186 119
rect -171 99 -169 119
rect -149 99 -147 119
rect -132 99 -130 119
rect -115 116 -113 120
rect -99 116 -97 120
rect -56 94 -54 104
rect -11 94 -9 104
rect 35 99 37 119
rect 52 99 54 119
rect 74 99 76 119
rect 91 99 93 119
rect 108 116 110 120
rect 124 116 126 120
rect 196 102 206 104
rect 232 98 234 108
rect 262 106 264 116
rect 298 102 308 104
rect 334 98 336 108
rect 364 106 366 116
rect 399 89 401 99
rect 444 89 446 99
rect 490 94 492 114
rect 507 94 509 114
rect 529 94 531 114
rect 546 94 548 114
rect 563 111 565 115
rect 579 111 581 115
rect -279 0 -277 10
rect -234 0 -232 10
rect -188 5 -186 25
rect -171 5 -169 25
rect -149 5 -147 25
rect -132 5 -130 25
rect -115 22 -113 26
rect -99 22 -97 26
rect 13 9 15 19
rect 43 17 45 27
rect 71 21 81 23
rect 197 30 207 32
rect 233 26 235 36
rect 263 34 265 44
rect 298 30 308 32
rect 334 26 336 36
rect 364 34 366 44
rect 19 -21 39 -19
rect 106 -27 108 -7
rect 122 -27 124 -7
rect 166 -17 168 -7
rect 409 -7 411 3
rect 454 -7 456 3
rect 500 -2 502 18
rect 517 -2 519 18
rect 539 -2 541 18
rect 556 -2 558 18
rect 573 15 575 19
rect 589 15 591 19
rect 143 -31 145 -21
rect 19 -37 39 -35
rect -279 -94 -277 -84
rect -234 -94 -232 -84
rect 29 -62 39 -60
rect -188 -89 -186 -69
rect -171 -89 -169 -69
rect -149 -89 -147 -69
rect -132 -89 -130 -69
rect -115 -72 -113 -68
rect -99 -72 -97 -68
rect 104 -108 106 -88
rect 120 -108 122 -88
rect 148 -98 150 -88
rect 190 -106 192 -86
rect 206 -106 208 -86
rect 250 -96 252 -86
rect 227 -110 229 -100
rect 284 -106 286 -86
rect 300 -106 302 -86
rect 344 -96 346 -86
rect 321 -110 323 -100
rect 378 -106 380 -86
rect 394 -106 396 -86
rect 438 -96 440 -86
rect 462 -98 464 -88
rect 507 -98 509 -88
rect 553 -93 555 -73
rect 570 -93 572 -73
rect 592 -93 594 -73
rect 609 -93 611 -73
rect 626 -76 628 -72
rect 642 -76 644 -72
rect 415 -110 417 -100
rect -6 -132 -4 -122
rect 24 -124 26 -114
rect 52 -120 62 -118
rect 448 -121 450 -111
rect -279 -187 -277 -177
rect -234 -187 -232 -177
rect 493 -121 495 -111
rect 539 -136 541 -116
rect 556 -136 558 -116
rect 578 -136 580 -116
rect 595 -136 597 -116
rect -188 -182 -186 -162
rect -171 -182 -169 -162
rect -149 -182 -147 -162
rect -132 -182 -130 -162
rect -115 -165 -113 -161
rect -99 -165 -97 -161
rect 0 -162 20 -160
rect 0 -178 20 -176
rect 328 -158 338 -156
rect 10 -203 20 -201
rect 104 -217 106 -177
rect 123 -217 125 -177
rect 142 -217 144 -177
rect 161 -217 163 -177
rect 177 -184 179 -174
rect 215 -192 217 -172
rect 231 -192 233 -172
rect 260 -182 262 -172
rect 612 -137 614 -133
rect 628 -137 630 -133
rect 328 -180 338 -178
rect 328 -200 338 -198
rect 509 -210 519 -208
rect -279 -281 -277 -271
rect -234 -281 -232 -271
rect -188 -276 -186 -256
rect -171 -276 -169 -256
rect -149 -276 -147 -256
rect -132 -276 -130 -256
rect -115 -259 -113 -255
rect -99 -259 -97 -255
rect -23 -273 -21 -263
rect 7 -265 9 -255
rect 328 -236 338 -234
rect 509 -255 519 -253
rect 35 -261 45 -259
rect -17 -303 3 -301
rect 112 -316 114 -276
rect 131 -316 133 -276
rect 150 -316 152 -276
rect 169 -316 171 -276
rect 185 -283 187 -273
rect 215 -286 217 -256
rect 231 -286 233 -256
rect 254 -286 256 -256
rect 279 -266 281 -256
rect 328 -257 338 -255
rect 328 -278 338 -276
rect 328 -299 338 -297
rect 494 -301 514 -299
rect -17 -319 3 -317
rect -279 -375 -277 -365
rect -234 -375 -232 -365
rect 494 -318 514 -316
rect -7 -344 3 -342
rect -188 -370 -186 -350
rect -171 -370 -169 -350
rect -149 -370 -147 -350
rect -132 -370 -130 -350
rect -115 -353 -113 -349
rect -99 -353 -97 -349
rect 494 -340 514 -338
rect 330 -344 340 -342
rect -41 -414 -39 -404
rect -11 -406 -9 -396
rect 17 -402 27 -400
rect 116 -405 118 -375
rect 132 -405 134 -375
rect 155 -405 157 -375
rect 180 -385 182 -375
rect 215 -380 217 -350
rect 231 -380 233 -350
rect 256 -380 258 -350
rect 284 -360 286 -350
rect 494 -357 514 -355
rect 330 -366 340 -364
rect 493 -374 497 -372
rect 330 -388 340 -386
rect 493 -390 497 -388
rect -279 -469 -277 -459
rect -234 -469 -232 -459
rect 330 -410 340 -408
rect -188 -464 -186 -444
rect -171 -464 -169 -444
rect -149 -464 -147 -444
rect -132 -464 -130 -444
rect -115 -447 -113 -443
rect -99 -447 -97 -443
rect -35 -444 -15 -442
rect 330 -431 340 -429
rect -35 -460 -15 -458
rect 215 -464 217 -444
rect 231 -464 233 -444
rect 256 -454 258 -444
rect -25 -485 -15 -483
rect 109 -489 111 -469
rect 125 -489 127 -469
rect 150 -479 152 -469
<< ptransistor >>
rect -279 120 -277 160
rect -257 120 -255 160
rect -234 120 -232 160
rect -212 120 -210 160
rect -179 143 -177 163
rect -140 143 -138 163
rect -115 141 -113 161
rect -99 141 -97 161
rect -56 120 -54 160
rect -34 120 -32 160
rect -11 120 -9 160
rect 11 120 13 160
rect 44 143 46 163
rect 83 143 85 163
rect 108 141 110 161
rect 124 141 126 161
rect 399 115 401 155
rect 421 115 423 155
rect 444 115 446 155
rect 466 115 468 155
rect 499 138 501 158
rect 538 138 540 158
rect 563 136 565 156
rect 579 136 581 156
rect 196 76 216 78
rect -279 26 -277 66
rect -257 26 -255 66
rect -234 26 -232 66
rect -212 26 -210 66
rect -179 49 -177 69
rect -140 49 -138 69
rect -115 47 -113 67
rect -99 47 -97 67
rect 232 63 234 83
rect 262 70 264 90
rect 298 76 318 78
rect 334 63 336 83
rect 364 70 366 90
rect 13 35 15 55
rect 43 42 45 62
rect 61 47 81 49
rect 106 9 108 49
rect 122 9 124 49
rect 143 9 145 49
rect 166 9 168 29
rect 55 -21 75 -19
rect -279 -68 -277 -28
rect -257 -68 -255 -28
rect -234 -68 -232 -28
rect -212 -68 -210 -28
rect -179 -45 -177 -25
rect -140 -45 -138 -25
rect 197 4 217 6
rect 233 -9 235 11
rect 263 -2 265 18
rect 409 19 411 59
rect 431 19 433 59
rect 454 19 456 59
rect 476 19 478 59
rect 509 42 511 62
rect 548 42 550 62
rect 573 40 575 60
rect 589 40 591 60
rect 298 4 318 6
rect 334 -9 336 11
rect 364 -2 366 18
rect -115 -47 -113 -27
rect -99 -47 -97 -27
rect 55 -37 75 -35
rect 55 -62 75 -60
rect 104 -72 106 -52
rect 120 -72 122 -52
rect 148 -72 150 -52
rect 190 -70 192 -30
rect 206 -70 208 -30
rect 227 -70 229 -30
rect 250 -70 252 -50
rect 284 -70 286 -30
rect 300 -70 302 -30
rect 321 -70 323 -30
rect 344 -70 346 -50
rect 378 -70 380 -30
rect 394 -70 396 -30
rect 415 -70 417 -30
rect 438 -70 440 -50
rect -6 -106 -4 -86
rect 24 -99 26 -79
rect 42 -94 62 -92
rect -279 -161 -277 -121
rect -257 -161 -255 -121
rect -234 -161 -232 -121
rect -212 -161 -210 -121
rect -179 -138 -177 -118
rect -140 -138 -138 -118
rect -115 -140 -113 -120
rect -99 -140 -97 -120
rect 462 -72 464 -32
rect 484 -72 486 -32
rect 507 -72 509 -32
rect 529 -72 531 -32
rect 562 -49 564 -29
rect 601 -49 603 -29
rect 626 -51 628 -31
rect 642 -51 644 -31
rect 104 -160 106 -140
rect 123 -160 125 -140
rect 142 -160 144 -140
rect 161 -160 163 -140
rect 177 -160 179 -140
rect 215 -156 217 -136
rect 231 -156 233 -136
rect 260 -156 262 -136
rect 36 -162 56 -160
rect 36 -178 56 -176
rect 354 -158 374 -156
rect 36 -203 56 -201
rect -279 -255 -277 -215
rect -257 -255 -255 -215
rect -234 -255 -232 -215
rect -212 -255 -210 -215
rect -179 -232 -177 -212
rect -140 -232 -138 -212
rect -115 -234 -113 -214
rect -99 -234 -97 -214
rect 448 -177 450 -137
rect 470 -177 472 -137
rect 493 -177 495 -137
rect 515 -177 517 -137
rect 354 -180 394 -178
rect 548 -180 550 -160
rect 587 -180 589 -160
rect 612 -178 614 -158
rect 628 -178 630 -158
rect 354 -200 394 -198
rect 453 -210 493 -208
rect -23 -247 -21 -227
rect 7 -240 9 -220
rect 25 -235 45 -233
rect 112 -259 114 -239
rect 131 -259 133 -239
rect 150 -259 152 -239
rect 169 -259 171 -239
rect 185 -259 187 -239
rect 215 -240 217 -220
rect 231 -240 233 -220
rect 254 -240 256 -220
rect 279 -240 281 -220
rect 453 -232 493 -230
rect 354 -236 374 -234
rect 453 -255 493 -253
rect 19 -303 39 -301
rect -279 -349 -277 -309
rect -257 -349 -255 -309
rect -234 -349 -232 -309
rect -212 -349 -210 -309
rect -179 -326 -177 -306
rect -140 -326 -138 -306
rect -115 -328 -113 -308
rect -99 -328 -97 -308
rect 354 -257 414 -255
rect 354 -278 414 -276
rect 453 -277 493 -275
rect 354 -299 414 -297
rect 450 -310 470 -308
rect 19 -319 39 -317
rect 215 -334 217 -314
rect 231 -334 233 -314
rect 256 -334 258 -314
rect 284 -334 286 -314
rect 19 -344 39 -342
rect 116 -359 118 -339
rect 132 -359 134 -339
rect 155 -359 157 -339
rect 180 -359 182 -339
rect 356 -344 376 -342
rect 450 -349 470 -347
rect -41 -388 -39 -368
rect -11 -381 -9 -361
rect 7 -376 27 -374
rect -279 -443 -277 -403
rect -257 -443 -255 -403
rect -234 -443 -232 -403
rect -212 -443 -210 -403
rect -179 -420 -177 -400
rect -140 -420 -138 -400
rect -115 -422 -113 -402
rect -99 -422 -97 -402
rect 356 -366 436 -364
rect 452 -374 472 -372
rect 356 -388 436 -386
rect 452 -390 472 -388
rect 215 -428 217 -408
rect 231 -428 233 -408
rect 256 -428 258 -408
rect 356 -410 436 -408
rect 1 -444 21 -442
rect 109 -453 111 -433
rect 125 -453 127 -433
rect 150 -453 152 -433
rect 356 -431 436 -429
rect 1 -460 21 -458
rect 1 -485 21 -483
<< ndiffusion >>
rect -280 94 -279 104
rect -277 94 -276 104
rect -235 94 -234 104
rect -232 94 -231 104
rect -189 99 -188 119
rect -186 99 -185 119
rect -172 99 -171 119
rect -169 99 -168 119
rect -150 99 -149 119
rect -147 99 -146 119
rect -133 99 -132 119
rect -130 99 -129 119
rect -116 116 -115 120
rect -113 116 -112 120
rect -100 116 -99 120
rect -97 116 -96 120
rect -57 94 -56 104
rect -54 94 -53 104
rect -12 94 -11 104
rect -9 94 -8 104
rect 34 99 35 119
rect 37 99 38 119
rect 51 99 52 119
rect 54 99 55 119
rect 73 99 74 119
rect 76 99 77 119
rect 90 99 91 119
rect 93 99 94 119
rect 107 116 108 120
rect 110 116 111 120
rect 123 116 124 120
rect 126 116 127 120
rect 196 104 206 105
rect 196 101 206 102
rect 231 98 232 108
rect 234 98 235 108
rect 261 106 262 116
rect 264 106 265 116
rect 298 104 308 105
rect 298 101 308 102
rect 333 98 334 108
rect 336 98 337 108
rect 363 106 364 116
rect 366 106 367 116
rect 398 89 399 99
rect 401 89 402 99
rect 443 89 444 99
rect 446 89 447 99
rect 489 94 490 114
rect 492 94 493 114
rect 506 94 507 114
rect 509 94 510 114
rect 528 94 529 114
rect 531 94 532 114
rect 545 94 546 114
rect 548 94 549 114
rect 562 111 563 115
rect 565 111 566 115
rect 578 111 579 115
rect 581 111 582 115
rect -280 0 -279 10
rect -277 0 -276 10
rect -235 0 -234 10
rect -232 0 -231 10
rect -189 5 -188 25
rect -186 5 -185 25
rect -172 5 -171 25
rect -169 5 -168 25
rect -150 5 -149 25
rect -147 5 -146 25
rect -133 5 -132 25
rect -130 5 -129 25
rect -116 22 -115 26
rect -113 22 -112 26
rect -100 22 -99 26
rect -97 22 -96 26
rect 12 9 13 19
rect 15 9 16 19
rect 42 17 43 27
rect 45 17 46 27
rect 71 23 81 24
rect 71 20 81 21
rect 197 32 207 33
rect 197 29 207 30
rect 232 26 233 36
rect 235 26 236 36
rect 262 34 263 44
rect 265 34 266 44
rect 298 32 308 33
rect 298 29 308 30
rect 333 26 334 36
rect 336 26 337 36
rect 363 34 364 44
rect 366 34 367 44
rect 19 -19 39 -18
rect 19 -22 39 -21
rect 105 -27 106 -7
rect 108 -27 109 -7
rect 121 -27 122 -7
rect 124 -27 125 -7
rect 165 -17 166 -7
rect 168 -17 169 -7
rect 408 -7 409 3
rect 411 -7 412 3
rect 453 -7 454 3
rect 456 -7 457 3
rect 499 -2 500 18
rect 502 -2 503 18
rect 516 -2 517 18
rect 519 -2 520 18
rect 538 -2 539 18
rect 541 -2 542 18
rect 555 -2 556 18
rect 558 -2 559 18
rect 572 15 573 19
rect 575 15 576 19
rect 588 15 589 19
rect 591 15 592 19
rect 19 -35 39 -34
rect 142 -31 143 -21
rect 145 -31 146 -21
rect 19 -38 39 -37
rect -280 -94 -279 -84
rect -277 -94 -276 -84
rect -235 -94 -234 -84
rect -232 -94 -231 -84
rect 29 -60 39 -59
rect 29 -63 39 -62
rect -189 -89 -188 -69
rect -186 -89 -185 -69
rect -172 -89 -171 -69
rect -169 -89 -168 -69
rect -150 -89 -149 -69
rect -147 -89 -146 -69
rect -133 -89 -132 -69
rect -130 -89 -129 -69
rect -116 -72 -115 -68
rect -113 -72 -112 -68
rect -100 -72 -99 -68
rect -97 -72 -96 -68
rect 103 -108 104 -88
rect 106 -108 107 -88
rect 119 -108 120 -88
rect 122 -108 123 -88
rect 147 -98 148 -88
rect 150 -98 151 -88
rect 189 -106 190 -86
rect 192 -106 193 -86
rect 205 -106 206 -86
rect 208 -106 209 -86
rect 249 -96 250 -86
rect 252 -96 253 -86
rect 226 -110 227 -100
rect 229 -110 230 -100
rect 283 -106 284 -86
rect 286 -106 287 -86
rect 299 -106 300 -86
rect 302 -106 303 -86
rect 343 -96 344 -86
rect 346 -96 347 -86
rect 320 -110 321 -100
rect 323 -110 324 -100
rect 377 -106 378 -86
rect 380 -106 381 -86
rect 393 -106 394 -86
rect 396 -106 397 -86
rect 437 -96 438 -86
rect 440 -96 441 -86
rect 461 -98 462 -88
rect 464 -98 465 -88
rect 506 -98 507 -88
rect 509 -98 510 -88
rect 552 -93 553 -73
rect 555 -93 556 -73
rect 569 -93 570 -73
rect 572 -93 573 -73
rect 591 -93 592 -73
rect 594 -93 595 -73
rect 608 -93 609 -73
rect 611 -93 612 -73
rect 625 -76 626 -72
rect 628 -76 629 -72
rect 641 -76 642 -72
rect 644 -76 645 -72
rect 414 -110 415 -100
rect 417 -110 418 -100
rect -7 -132 -6 -122
rect -4 -132 -3 -122
rect 23 -124 24 -114
rect 26 -124 27 -114
rect 52 -118 62 -117
rect 52 -121 62 -120
rect 447 -121 448 -111
rect 450 -121 451 -111
rect -280 -187 -279 -177
rect -277 -187 -276 -177
rect -235 -187 -234 -177
rect -232 -187 -231 -177
rect 0 -160 20 -159
rect 492 -121 493 -111
rect 495 -121 496 -111
rect 538 -136 539 -116
rect 541 -136 542 -116
rect 555 -136 556 -116
rect 558 -136 559 -116
rect 577 -136 578 -116
rect 580 -136 581 -116
rect 594 -136 595 -116
rect 597 -136 598 -116
rect 328 -156 338 -155
rect -189 -182 -188 -162
rect -186 -182 -185 -162
rect -172 -182 -171 -162
rect -169 -182 -168 -162
rect -150 -182 -149 -162
rect -147 -182 -146 -162
rect -133 -182 -132 -162
rect -130 -182 -129 -162
rect -116 -165 -115 -161
rect -113 -165 -112 -161
rect -100 -165 -99 -161
rect -97 -165 -96 -161
rect 0 -163 20 -162
rect 0 -176 20 -175
rect 328 -159 338 -158
rect 0 -179 20 -178
rect 10 -201 20 -200
rect 10 -204 20 -203
rect 103 -217 104 -177
rect 106 -217 107 -177
rect 122 -217 123 -177
rect 125 -217 126 -177
rect 141 -217 142 -177
rect 144 -217 145 -177
rect 160 -217 161 -177
rect 163 -217 164 -177
rect 176 -184 177 -174
rect 179 -184 180 -174
rect 214 -192 215 -172
rect 217 -192 218 -172
rect 230 -192 231 -172
rect 233 -192 234 -172
rect 259 -182 260 -172
rect 262 -182 263 -172
rect 328 -178 338 -177
rect 611 -137 612 -133
rect 614 -137 615 -133
rect 627 -137 628 -133
rect 630 -137 631 -133
rect 328 -181 338 -180
rect 328 -198 338 -197
rect 328 -201 338 -200
rect 509 -208 519 -207
rect 509 -211 519 -210
rect -280 -281 -279 -271
rect -277 -281 -276 -271
rect -235 -281 -234 -271
rect -232 -281 -231 -271
rect -189 -276 -188 -256
rect -186 -276 -185 -256
rect -172 -276 -171 -256
rect -169 -276 -168 -256
rect -150 -276 -149 -256
rect -147 -276 -146 -256
rect -133 -276 -132 -256
rect -130 -276 -129 -256
rect -116 -259 -115 -255
rect -113 -259 -112 -255
rect -100 -259 -99 -255
rect -97 -259 -96 -255
rect -24 -273 -23 -263
rect -21 -273 -20 -263
rect 6 -265 7 -255
rect 9 -265 10 -255
rect 35 -259 45 -258
rect 328 -234 338 -233
rect 328 -237 338 -236
rect 328 -255 338 -254
rect 509 -253 519 -252
rect 35 -262 45 -261
rect -17 -301 3 -300
rect -17 -304 3 -303
rect -17 -317 3 -316
rect 111 -316 112 -276
rect 114 -316 115 -276
rect 130 -316 131 -276
rect 133 -316 134 -276
rect 149 -316 150 -276
rect 152 -316 153 -276
rect 168 -316 169 -276
rect 171 -316 172 -276
rect 184 -283 185 -273
rect 187 -283 188 -273
rect 214 -286 215 -256
rect 217 -286 218 -256
rect 230 -286 231 -256
rect 233 -286 234 -256
rect 253 -286 254 -256
rect 256 -286 257 -256
rect 278 -266 279 -256
rect 281 -266 282 -256
rect 328 -258 338 -257
rect 509 -256 519 -255
rect 328 -276 338 -275
rect 328 -279 338 -278
rect 328 -297 338 -296
rect 494 -299 514 -298
rect 328 -300 338 -299
rect 494 -302 514 -301
rect -17 -320 3 -319
rect -280 -375 -279 -365
rect -277 -375 -276 -365
rect -235 -375 -234 -365
rect -232 -375 -231 -365
rect 494 -316 514 -315
rect 494 -319 514 -318
rect -7 -342 3 -341
rect -7 -345 3 -344
rect -189 -370 -188 -350
rect -186 -370 -185 -350
rect -172 -370 -171 -350
rect -169 -370 -168 -350
rect -150 -370 -149 -350
rect -147 -370 -146 -350
rect -133 -370 -132 -350
rect -130 -370 -129 -350
rect -116 -353 -115 -349
rect -113 -353 -112 -349
rect -100 -353 -99 -349
rect -97 -353 -96 -349
rect 330 -342 340 -341
rect 494 -338 514 -337
rect 494 -341 514 -340
rect 330 -345 340 -344
rect -42 -414 -41 -404
rect -39 -414 -38 -404
rect -12 -406 -11 -396
rect -9 -406 -8 -396
rect 17 -400 27 -399
rect 17 -403 27 -402
rect 115 -405 116 -375
rect 118 -405 119 -375
rect 131 -405 132 -375
rect 134 -405 135 -375
rect 154 -405 155 -375
rect 157 -405 158 -375
rect 179 -385 180 -375
rect 182 -385 183 -375
rect 214 -380 215 -350
rect 217 -380 218 -350
rect 230 -380 231 -350
rect 233 -380 234 -350
rect 255 -380 256 -350
rect 258 -380 259 -350
rect 283 -360 284 -350
rect 286 -360 287 -350
rect 494 -355 514 -354
rect 494 -358 514 -357
rect 330 -364 340 -363
rect 330 -367 340 -366
rect 493 -372 497 -371
rect 493 -375 497 -374
rect 330 -386 340 -385
rect 493 -388 497 -387
rect 330 -389 340 -388
rect 493 -391 497 -390
rect 330 -408 340 -407
rect -280 -469 -279 -459
rect -277 -469 -276 -459
rect -235 -469 -234 -459
rect -232 -469 -231 -459
rect 330 -411 340 -410
rect -35 -442 -15 -441
rect -189 -464 -188 -444
rect -186 -464 -185 -444
rect -172 -464 -171 -444
rect -169 -464 -168 -444
rect -150 -464 -149 -444
rect -147 -464 -146 -444
rect -133 -464 -132 -444
rect -130 -464 -129 -444
rect -116 -447 -115 -443
rect -113 -447 -112 -443
rect -100 -447 -99 -443
rect -97 -447 -96 -443
rect -35 -445 -15 -444
rect 330 -429 340 -428
rect 330 -432 340 -431
rect -35 -458 -15 -457
rect -35 -461 -15 -460
rect 214 -464 215 -444
rect 217 -464 218 -444
rect 230 -464 231 -444
rect 233 -464 234 -444
rect 255 -454 256 -444
rect 258 -454 259 -444
rect -25 -483 -15 -482
rect -25 -486 -15 -485
rect 108 -489 109 -469
rect 111 -489 112 -469
rect 124 -489 125 -469
rect 127 -489 128 -469
rect 149 -479 150 -469
rect 152 -479 153 -469
<< pdiffusion >>
rect -280 120 -279 160
rect -277 120 -276 160
rect -258 120 -257 160
rect -255 120 -254 160
rect -235 120 -234 160
rect -232 120 -231 160
rect -213 120 -212 160
rect -210 120 -209 160
rect -180 143 -179 163
rect -177 143 -176 163
rect -141 143 -140 163
rect -138 143 -137 163
rect -116 141 -115 161
rect -113 141 -112 161
rect -100 141 -99 161
rect -97 141 -96 161
rect -57 120 -56 160
rect -54 120 -53 160
rect -35 120 -34 160
rect -32 120 -31 160
rect -12 120 -11 160
rect -9 120 -8 160
rect 10 120 11 160
rect 13 120 14 160
rect 43 143 44 163
rect 46 143 47 163
rect 82 143 83 163
rect 85 143 86 163
rect 107 141 108 161
rect 110 141 111 161
rect 123 141 124 161
rect 126 141 127 161
rect 398 115 399 155
rect 401 115 402 155
rect 420 115 421 155
rect 423 115 424 155
rect 443 115 444 155
rect 446 115 447 155
rect 465 115 466 155
rect 468 115 469 155
rect 498 138 499 158
rect 501 138 502 158
rect 537 138 538 158
rect 540 138 541 158
rect 562 136 563 156
rect 565 136 566 156
rect 578 136 579 156
rect 581 136 582 156
rect 196 78 216 79
rect 196 75 216 76
rect -280 26 -279 66
rect -277 26 -276 66
rect -258 26 -257 66
rect -255 26 -254 66
rect -235 26 -234 66
rect -232 26 -231 66
rect -213 26 -212 66
rect -210 26 -209 66
rect -180 49 -179 69
rect -177 49 -176 69
rect -141 49 -140 69
rect -138 49 -137 69
rect -116 47 -115 67
rect -113 47 -112 67
rect -100 47 -99 67
rect -97 47 -96 67
rect 231 63 232 83
rect 234 63 235 83
rect 261 70 262 90
rect 264 70 265 90
rect 298 78 318 79
rect 298 75 318 76
rect 333 63 334 83
rect 336 63 337 83
rect 363 70 364 90
rect 366 70 367 90
rect 12 35 13 55
rect 15 35 16 55
rect 42 42 43 62
rect 45 42 46 62
rect 61 49 81 50
rect 61 46 81 47
rect 105 9 106 49
rect 108 9 109 49
rect 121 9 122 49
rect 124 9 125 49
rect 142 9 143 49
rect 145 9 146 49
rect 165 9 166 29
rect 168 9 169 29
rect 55 -19 75 -18
rect -280 -68 -279 -28
rect -277 -68 -276 -28
rect -258 -68 -257 -28
rect -255 -68 -254 -28
rect -235 -68 -234 -28
rect -232 -68 -231 -28
rect -213 -68 -212 -28
rect -210 -68 -209 -28
rect -180 -45 -179 -25
rect -177 -45 -176 -25
rect -141 -45 -140 -25
rect -138 -45 -137 -25
rect 55 -22 75 -21
rect 197 6 217 7
rect 197 3 217 4
rect 232 -9 233 11
rect 235 -9 236 11
rect 262 -2 263 18
rect 265 -2 266 18
rect 408 19 409 59
rect 411 19 412 59
rect 430 19 431 59
rect 433 19 434 59
rect 453 19 454 59
rect 456 19 457 59
rect 475 19 476 59
rect 478 19 479 59
rect 508 42 509 62
rect 511 42 512 62
rect 547 42 548 62
rect 550 42 551 62
rect 572 40 573 60
rect 575 40 576 60
rect 588 40 589 60
rect 591 40 592 60
rect 298 6 318 7
rect 298 3 318 4
rect 333 -9 334 11
rect 336 -9 337 11
rect 363 -2 364 18
rect 366 -2 367 18
rect -116 -47 -115 -27
rect -113 -47 -112 -27
rect -100 -47 -99 -27
rect -97 -47 -96 -27
rect 55 -35 75 -34
rect 55 -38 75 -37
rect 55 -60 75 -59
rect 55 -63 75 -62
rect 103 -72 104 -52
rect 106 -72 107 -52
rect 119 -72 120 -52
rect 122 -72 123 -52
rect 147 -72 148 -52
rect 150 -72 151 -52
rect 189 -70 190 -30
rect 192 -70 193 -30
rect 205 -70 206 -30
rect 208 -70 209 -30
rect 226 -70 227 -30
rect 229 -70 230 -30
rect 249 -70 250 -50
rect 252 -70 253 -50
rect 283 -70 284 -30
rect 286 -70 287 -30
rect 299 -70 300 -30
rect 302 -70 303 -30
rect 320 -70 321 -30
rect 323 -70 324 -30
rect 343 -70 344 -50
rect 346 -70 347 -50
rect 377 -70 378 -30
rect 380 -70 381 -30
rect 393 -70 394 -30
rect 396 -70 397 -30
rect 414 -70 415 -30
rect 417 -70 418 -30
rect 437 -70 438 -50
rect 440 -70 441 -50
rect -7 -106 -6 -86
rect -4 -106 -3 -86
rect 23 -99 24 -79
rect 26 -99 27 -79
rect 42 -92 62 -91
rect 42 -95 62 -94
rect -280 -161 -279 -121
rect -277 -161 -276 -121
rect -258 -161 -257 -121
rect -255 -161 -254 -121
rect -235 -161 -234 -121
rect -232 -161 -231 -121
rect -213 -161 -212 -121
rect -210 -161 -209 -121
rect -180 -138 -179 -118
rect -177 -138 -176 -118
rect -141 -138 -140 -118
rect -138 -138 -137 -118
rect -116 -140 -115 -120
rect -113 -140 -112 -120
rect -100 -140 -99 -120
rect -97 -140 -96 -120
rect 461 -72 462 -32
rect 464 -72 465 -32
rect 483 -72 484 -32
rect 486 -72 487 -32
rect 506 -72 507 -32
rect 509 -72 510 -32
rect 528 -72 529 -32
rect 531 -72 532 -32
rect 561 -49 562 -29
rect 564 -49 565 -29
rect 600 -49 601 -29
rect 603 -49 604 -29
rect 625 -51 626 -31
rect 628 -51 629 -31
rect 641 -51 642 -31
rect 644 -51 645 -31
rect 36 -160 56 -159
rect 103 -160 104 -140
rect 106 -160 107 -140
rect 122 -160 123 -140
rect 125 -160 126 -140
rect 141 -160 142 -140
rect 144 -160 145 -140
rect 160 -160 161 -140
rect 163 -160 164 -140
rect 176 -160 177 -140
rect 179 -160 180 -140
rect 214 -156 215 -136
rect 217 -156 218 -136
rect 230 -156 231 -136
rect 233 -156 234 -136
rect 259 -156 260 -136
rect 262 -156 263 -136
rect 354 -156 374 -155
rect 36 -163 56 -162
rect 36 -176 56 -175
rect 354 -159 374 -158
rect 36 -179 56 -178
rect 36 -201 56 -200
rect 36 -204 56 -203
rect -280 -255 -279 -215
rect -277 -255 -276 -215
rect -258 -255 -257 -215
rect -255 -255 -254 -215
rect -235 -255 -234 -215
rect -232 -255 -231 -215
rect -213 -255 -212 -215
rect -210 -255 -209 -215
rect -180 -232 -179 -212
rect -177 -232 -176 -212
rect -141 -232 -140 -212
rect -138 -232 -137 -212
rect -116 -234 -115 -214
rect -113 -234 -112 -214
rect -100 -234 -99 -214
rect -97 -234 -96 -214
rect 447 -177 448 -137
rect 450 -177 451 -137
rect 469 -177 470 -137
rect 472 -177 473 -137
rect 492 -177 493 -137
rect 495 -177 496 -137
rect 514 -177 515 -137
rect 517 -177 518 -137
rect 354 -178 394 -177
rect 547 -180 548 -160
rect 550 -180 551 -160
rect 586 -180 587 -160
rect 589 -180 590 -160
rect 611 -178 612 -158
rect 614 -178 615 -158
rect 627 -178 628 -158
rect 630 -178 631 -158
rect 354 -181 394 -180
rect 354 -198 394 -197
rect 354 -201 394 -200
rect 453 -208 493 -207
rect 453 -211 493 -210
rect -24 -247 -23 -227
rect -21 -247 -20 -227
rect 6 -240 7 -220
rect 9 -240 10 -220
rect 25 -233 45 -232
rect 25 -236 45 -235
rect 111 -259 112 -239
rect 114 -259 115 -239
rect 130 -259 131 -239
rect 133 -259 134 -239
rect 149 -259 150 -239
rect 152 -259 153 -239
rect 168 -259 169 -239
rect 171 -259 172 -239
rect 184 -259 185 -239
rect 187 -259 188 -239
rect 214 -240 215 -220
rect 217 -240 218 -220
rect 230 -240 231 -220
rect 233 -240 234 -220
rect 253 -240 254 -220
rect 256 -240 257 -220
rect 278 -240 279 -220
rect 281 -240 282 -220
rect 453 -230 493 -229
rect 354 -234 374 -233
rect 453 -233 493 -232
rect 354 -237 374 -236
rect 453 -253 493 -252
rect 354 -255 414 -254
rect 19 -301 39 -300
rect -280 -349 -279 -309
rect -277 -349 -276 -309
rect -258 -349 -257 -309
rect -255 -349 -254 -309
rect -235 -349 -234 -309
rect -232 -349 -231 -309
rect -213 -349 -212 -309
rect -210 -349 -209 -309
rect -180 -326 -179 -306
rect -177 -326 -176 -306
rect -141 -326 -140 -306
rect -138 -326 -137 -306
rect 19 -304 39 -303
rect -116 -328 -115 -308
rect -113 -328 -112 -308
rect -100 -328 -99 -308
rect -97 -328 -96 -308
rect 453 -256 493 -255
rect 354 -258 414 -257
rect 453 -275 493 -274
rect 354 -276 414 -275
rect 453 -278 493 -277
rect 354 -279 414 -278
rect 354 -297 414 -296
rect 354 -300 414 -299
rect 450 -308 470 -307
rect 450 -311 470 -310
rect 19 -317 39 -316
rect 19 -320 39 -319
rect 214 -334 215 -314
rect 217 -334 218 -314
rect 230 -334 231 -314
rect 233 -334 234 -314
rect 255 -334 256 -314
rect 258 -334 259 -314
rect 283 -334 284 -314
rect 286 -334 287 -314
rect 19 -342 39 -341
rect 19 -345 39 -344
rect 115 -359 116 -339
rect 118 -359 119 -339
rect 131 -359 132 -339
rect 134 -359 135 -339
rect 154 -359 155 -339
rect 157 -359 158 -339
rect 179 -359 180 -339
rect 182 -359 183 -339
rect 356 -342 376 -341
rect 356 -345 376 -344
rect 450 -347 470 -346
rect 450 -350 470 -349
rect -42 -388 -41 -368
rect -39 -388 -38 -368
rect -12 -381 -11 -361
rect -9 -381 -8 -361
rect 7 -374 27 -373
rect 7 -377 27 -376
rect -280 -443 -279 -403
rect -277 -443 -276 -403
rect -258 -443 -257 -403
rect -255 -443 -254 -403
rect -235 -443 -234 -403
rect -232 -443 -231 -403
rect -213 -443 -212 -403
rect -210 -443 -209 -403
rect -180 -420 -179 -400
rect -177 -420 -176 -400
rect -141 -420 -140 -400
rect -138 -420 -137 -400
rect -116 -422 -115 -402
rect -113 -422 -112 -402
rect -100 -422 -99 -402
rect -97 -422 -96 -402
rect 356 -364 436 -363
rect 356 -367 436 -366
rect 452 -372 472 -371
rect 452 -375 472 -374
rect 356 -386 436 -385
rect 452 -388 472 -387
rect 356 -389 436 -388
rect 452 -391 472 -390
rect 356 -408 436 -407
rect 214 -428 215 -408
rect 217 -428 218 -408
rect 230 -428 231 -408
rect 233 -428 234 -408
rect 255 -428 256 -408
rect 258 -428 259 -408
rect 356 -411 436 -410
rect 1 -442 21 -441
rect 1 -445 21 -444
rect 108 -453 109 -433
rect 111 -453 112 -433
rect 124 -453 125 -433
rect 127 -453 128 -433
rect 149 -453 150 -433
rect 152 -453 153 -433
rect 356 -429 436 -428
rect 356 -432 436 -431
rect 1 -458 21 -457
rect 1 -461 21 -460
rect 1 -483 21 -482
rect 1 -486 21 -485
<< ndcontact >>
rect -284 94 -280 104
rect -276 94 -271 104
rect -239 94 -235 104
rect -231 94 -226 104
rect -193 99 -189 119
rect -185 99 -180 119
rect -176 99 -172 119
rect -168 99 -163 119
rect -154 99 -150 119
rect -146 99 -141 119
rect -137 99 -133 119
rect -129 99 -124 119
rect -120 116 -116 120
rect -112 116 -108 120
rect -104 116 -100 120
rect -96 116 -92 120
rect -61 94 -57 104
rect -53 94 -48 104
rect -16 94 -12 104
rect -8 94 -3 104
rect 30 99 34 119
rect 38 99 43 119
rect 47 99 51 119
rect 55 99 60 119
rect 69 99 73 119
rect 77 99 82 119
rect 86 99 90 119
rect 94 99 99 119
rect 103 116 107 120
rect 111 116 115 120
rect 119 116 123 120
rect 127 116 131 120
rect 196 105 206 109
rect 196 97 206 101
rect 227 98 231 108
rect 235 98 239 108
rect 257 106 261 116
rect 265 106 269 116
rect 298 105 308 109
rect 298 97 308 101
rect 329 98 333 108
rect 337 98 341 108
rect 359 106 363 116
rect 367 106 371 116
rect 394 89 398 99
rect 402 89 407 99
rect 439 89 443 99
rect 447 89 452 99
rect 485 94 489 114
rect 493 94 498 114
rect 502 94 506 114
rect 510 94 515 114
rect 524 94 528 114
rect 532 94 537 114
rect 541 94 545 114
rect 549 94 554 114
rect 558 111 562 115
rect 566 111 570 115
rect 574 111 578 115
rect 582 111 586 115
rect -284 0 -280 10
rect -276 0 -271 10
rect -239 0 -235 10
rect -231 0 -226 10
rect -193 5 -189 25
rect -185 5 -180 25
rect -176 5 -172 25
rect -168 5 -163 25
rect -154 5 -150 25
rect -146 5 -141 25
rect -137 5 -133 25
rect -129 5 -124 25
rect -120 22 -116 26
rect -112 22 -108 26
rect -104 22 -100 26
rect -96 22 -92 26
rect 8 9 12 19
rect 16 9 20 19
rect 38 17 42 27
rect 46 17 50 27
rect 71 24 81 28
rect 71 16 81 20
rect 197 33 207 37
rect 197 25 207 29
rect 228 26 232 36
rect 236 26 240 36
rect 258 34 262 44
rect 266 34 270 44
rect 298 33 308 37
rect 298 25 308 29
rect 329 26 333 36
rect 337 26 341 36
rect 359 34 363 44
rect 367 34 371 44
rect 19 -18 39 -14
rect 19 -26 39 -22
rect 101 -27 105 -7
rect 109 -27 113 -7
rect 117 -27 121 -7
rect 125 -27 129 -7
rect 161 -17 165 -7
rect 169 -17 173 -7
rect 404 -7 408 3
rect 412 -7 417 3
rect 449 -7 453 3
rect 457 -7 462 3
rect 495 -2 499 18
rect 503 -2 508 18
rect 512 -2 516 18
rect 520 -2 525 18
rect 534 -2 538 18
rect 542 -2 547 18
rect 551 -2 555 18
rect 559 -2 564 18
rect 568 15 572 19
rect 576 15 580 19
rect 584 15 588 19
rect 592 15 596 19
rect 19 -34 39 -30
rect 138 -31 142 -21
rect 146 -31 150 -21
rect 19 -42 39 -38
rect -284 -94 -280 -84
rect -276 -94 -271 -84
rect -239 -94 -235 -84
rect -231 -94 -226 -84
rect 29 -59 39 -55
rect 29 -67 39 -63
rect -193 -89 -189 -69
rect -185 -89 -180 -69
rect -176 -89 -172 -69
rect -168 -89 -163 -69
rect -154 -89 -150 -69
rect -146 -89 -141 -69
rect -137 -89 -133 -69
rect -129 -89 -124 -69
rect -120 -72 -116 -68
rect -112 -72 -108 -68
rect -104 -72 -100 -68
rect -96 -72 -92 -68
rect 99 -108 103 -88
rect 107 -108 111 -88
rect 115 -108 119 -88
rect 123 -108 127 -88
rect 143 -98 147 -88
rect 151 -98 155 -88
rect 185 -106 189 -86
rect 193 -106 197 -86
rect 201 -106 205 -86
rect 209 -106 213 -86
rect 245 -96 249 -86
rect 253 -96 257 -86
rect 222 -110 226 -100
rect 230 -110 234 -100
rect 279 -106 283 -86
rect 287 -106 291 -86
rect 295 -106 299 -86
rect 303 -106 307 -86
rect 339 -96 343 -86
rect 347 -96 351 -86
rect 316 -110 320 -100
rect 324 -110 328 -100
rect 373 -106 377 -86
rect 381 -106 385 -86
rect 389 -106 393 -86
rect 397 -106 401 -86
rect 433 -96 437 -86
rect 441 -96 445 -86
rect 457 -98 461 -88
rect 465 -98 470 -88
rect 502 -98 506 -88
rect 510 -98 515 -88
rect 548 -93 552 -73
rect 556 -93 561 -73
rect 565 -93 569 -73
rect 573 -93 578 -73
rect 587 -93 591 -73
rect 595 -93 600 -73
rect 604 -93 608 -73
rect 612 -93 617 -73
rect 621 -76 625 -72
rect 629 -76 633 -72
rect 637 -76 641 -72
rect 645 -76 649 -72
rect 410 -110 414 -100
rect 418 -110 422 -100
rect -11 -132 -7 -122
rect -3 -132 1 -122
rect 19 -124 23 -114
rect 27 -124 31 -114
rect 52 -117 62 -113
rect 443 -121 447 -111
rect 451 -121 456 -111
rect 52 -125 62 -121
rect -284 -187 -280 -177
rect -276 -187 -271 -177
rect -239 -187 -235 -177
rect -231 -187 -226 -177
rect 0 -159 20 -155
rect 488 -121 492 -111
rect 496 -121 501 -111
rect 534 -136 538 -116
rect 542 -136 547 -116
rect 551 -136 555 -116
rect 559 -136 564 -116
rect 573 -136 577 -116
rect 581 -136 586 -116
rect 590 -136 594 -116
rect 598 -136 603 -116
rect 328 -155 338 -151
rect -193 -182 -189 -162
rect -185 -182 -180 -162
rect -176 -182 -172 -162
rect -168 -182 -163 -162
rect -154 -182 -150 -162
rect -146 -182 -141 -162
rect -137 -182 -133 -162
rect -129 -182 -124 -162
rect -120 -165 -116 -161
rect -112 -165 -108 -161
rect -104 -165 -100 -161
rect -96 -165 -92 -161
rect 0 -167 20 -163
rect 0 -175 20 -171
rect 328 -163 338 -159
rect 0 -183 20 -179
rect 10 -200 20 -196
rect 10 -208 20 -204
rect 99 -217 103 -177
rect 107 -217 111 -177
rect 118 -217 122 -177
rect 126 -217 130 -177
rect 137 -217 141 -177
rect 145 -217 149 -177
rect 156 -217 160 -177
rect 164 -217 168 -177
rect 172 -184 176 -174
rect 180 -184 184 -174
rect 210 -192 214 -172
rect 218 -192 222 -172
rect 226 -192 230 -172
rect 234 -192 238 -172
rect 255 -182 259 -172
rect 263 -182 267 -172
rect 328 -177 338 -172
rect 607 -137 611 -133
rect 615 -137 619 -133
rect 623 -137 627 -133
rect 631 -137 635 -133
rect 328 -185 338 -181
rect 328 -197 338 -192
rect 328 -206 338 -201
rect 509 -207 519 -203
rect 509 -216 519 -211
rect -284 -281 -280 -271
rect -276 -281 -271 -271
rect -239 -281 -235 -271
rect -231 -281 -226 -271
rect -193 -276 -189 -256
rect -185 -276 -180 -256
rect -176 -276 -172 -256
rect -168 -276 -163 -256
rect -154 -276 -150 -256
rect -146 -276 -141 -256
rect -137 -276 -133 -256
rect -129 -276 -124 -256
rect -120 -259 -116 -255
rect -112 -259 -108 -255
rect -104 -259 -100 -255
rect -96 -259 -92 -255
rect -28 -273 -24 -263
rect -20 -273 -16 -263
rect 2 -265 6 -255
rect 10 -265 14 -255
rect 35 -258 45 -254
rect 328 -233 338 -229
rect 328 -241 338 -237
rect 328 -254 338 -249
rect 509 -252 519 -248
rect 35 -266 45 -262
rect -17 -300 3 -296
rect -17 -308 3 -304
rect -17 -316 3 -312
rect 107 -316 111 -276
rect 115 -316 119 -276
rect 126 -316 130 -276
rect 134 -316 138 -276
rect 145 -316 149 -276
rect 153 -316 157 -276
rect 164 -316 168 -276
rect 172 -316 176 -276
rect 180 -283 184 -273
rect 188 -283 192 -273
rect 210 -286 214 -256
rect 218 -286 222 -256
rect 226 -286 230 -256
rect 234 -286 238 -256
rect 249 -286 253 -256
rect 257 -286 261 -256
rect 274 -266 278 -256
rect 282 -266 286 -256
rect 328 -262 338 -258
rect 509 -261 519 -256
rect 328 -275 338 -270
rect 328 -284 338 -279
rect 328 -296 338 -291
rect 494 -298 514 -294
rect 328 -305 338 -300
rect 494 -307 514 -302
rect -17 -324 3 -320
rect -284 -375 -280 -365
rect -276 -375 -271 -365
rect -239 -375 -235 -365
rect -231 -375 -226 -365
rect 494 -315 514 -311
rect 494 -324 514 -319
rect -7 -341 3 -337
rect -7 -349 3 -345
rect -193 -370 -189 -350
rect -185 -370 -180 -350
rect -176 -370 -172 -350
rect -168 -370 -163 -350
rect -154 -370 -150 -350
rect -146 -370 -141 -350
rect -137 -370 -133 -350
rect -129 -370 -124 -350
rect -120 -353 -116 -349
rect -112 -353 -108 -349
rect -104 -353 -100 -349
rect -96 -353 -92 -349
rect 330 -341 340 -337
rect 494 -337 514 -333
rect 330 -349 340 -345
rect 494 -346 514 -341
rect -46 -414 -42 -404
rect -38 -414 -34 -404
rect -16 -406 -12 -396
rect -8 -406 -4 -396
rect 17 -399 27 -395
rect 17 -407 27 -403
rect 111 -405 115 -375
rect 119 -405 123 -375
rect 127 -405 131 -375
rect 135 -405 139 -375
rect 150 -405 154 -375
rect 158 -405 162 -375
rect 175 -385 179 -375
rect 183 -385 187 -375
rect 210 -380 214 -350
rect 218 -380 222 -350
rect 226 -380 230 -350
rect 234 -380 238 -350
rect 251 -380 255 -350
rect 259 -380 263 -350
rect 279 -360 283 -350
rect 287 -360 291 -350
rect 494 -354 514 -350
rect 330 -363 340 -358
rect 494 -363 514 -358
rect 330 -371 340 -367
rect 493 -371 497 -367
rect 493 -379 497 -375
rect 330 -385 340 -380
rect 493 -387 497 -383
rect 330 -394 340 -389
rect 493 -395 497 -391
rect 330 -407 340 -402
rect -284 -469 -280 -459
rect -276 -469 -271 -459
rect -239 -469 -235 -459
rect -231 -469 -226 -459
rect 330 -416 340 -411
rect 330 -428 340 -423
rect -35 -441 -15 -437
rect -193 -464 -189 -444
rect -185 -464 -180 -444
rect -176 -464 -172 -444
rect -168 -464 -163 -444
rect -154 -464 -150 -444
rect -146 -464 -141 -444
rect -137 -464 -133 -444
rect -129 -464 -124 -444
rect -120 -447 -116 -443
rect -112 -447 -108 -443
rect -104 -447 -100 -443
rect -96 -447 -92 -443
rect -35 -449 -15 -445
rect 330 -437 340 -432
rect -35 -457 -15 -453
rect -35 -465 -15 -461
rect 210 -464 214 -444
rect 218 -464 222 -444
rect 226 -464 230 -444
rect 234 -464 238 -444
rect 251 -454 255 -444
rect 259 -454 263 -444
rect -25 -482 -15 -478
rect -25 -490 -15 -486
rect 104 -489 108 -469
rect 112 -489 116 -469
rect 120 -489 124 -469
rect 128 -489 132 -469
rect 145 -479 149 -469
rect 153 -479 157 -469
<< pdcontact >>
rect -284 120 -280 160
rect -276 120 -272 160
rect -262 120 -258 160
rect -254 120 -250 160
rect -239 120 -235 160
rect -231 120 -227 160
rect -217 120 -213 160
rect -209 120 -205 160
rect -185 143 -180 163
rect -176 143 -172 163
rect -146 143 -141 163
rect -137 143 -133 163
rect -120 141 -116 161
rect -112 141 -108 161
rect -104 141 -100 161
rect -96 141 -92 161
rect -61 120 -57 160
rect -53 120 -49 160
rect -39 120 -35 160
rect -31 120 -27 160
rect -16 120 -12 160
rect -8 120 -4 160
rect 6 120 10 160
rect 14 120 18 160
rect 38 143 43 163
rect 47 143 51 163
rect 77 143 82 163
rect 86 143 90 163
rect 103 141 107 161
rect 111 141 115 161
rect 119 141 123 161
rect 127 141 131 161
rect 394 115 398 155
rect 402 115 406 155
rect 416 115 420 155
rect 424 115 428 155
rect 439 115 443 155
rect 447 115 451 155
rect 461 115 465 155
rect 469 115 473 155
rect 493 138 498 158
rect 502 138 506 158
rect 532 138 537 158
rect 541 138 545 158
rect 558 136 562 156
rect 566 136 570 156
rect 574 136 578 156
rect 582 136 586 156
rect 196 79 216 83
rect 196 71 216 75
rect -284 26 -280 66
rect -276 26 -272 66
rect -262 26 -258 66
rect -254 26 -250 66
rect -239 26 -235 66
rect -231 26 -227 66
rect -217 26 -213 66
rect -209 26 -205 66
rect -185 49 -180 69
rect -176 49 -172 69
rect -146 49 -141 69
rect -137 49 -133 69
rect -120 47 -116 67
rect -112 47 -108 67
rect -104 47 -100 67
rect -96 47 -92 67
rect 227 63 231 83
rect 235 63 239 83
rect 257 70 261 90
rect 265 70 269 90
rect 298 79 318 83
rect 298 71 318 75
rect 329 63 333 83
rect 337 63 341 83
rect 359 70 363 90
rect 367 70 371 90
rect 8 35 12 55
rect 16 35 20 55
rect 38 42 42 62
rect 46 42 50 62
rect 61 50 81 54
rect 61 42 81 46
rect 101 9 105 49
rect 109 9 113 49
rect 117 9 121 49
rect 125 9 129 49
rect 138 9 142 49
rect 146 9 150 49
rect 161 9 165 29
rect 169 9 173 29
rect 55 -18 75 -14
rect -284 -68 -280 -28
rect -276 -68 -272 -28
rect -262 -68 -258 -28
rect -254 -68 -250 -28
rect -239 -68 -235 -28
rect -231 -68 -227 -28
rect -217 -68 -213 -28
rect -209 -68 -205 -28
rect -185 -45 -180 -25
rect -176 -45 -172 -25
rect -146 -45 -141 -25
rect -137 -45 -133 -25
rect 55 -26 75 -22
rect 197 7 217 11
rect 197 -1 217 3
rect 228 -9 232 11
rect 236 -9 240 11
rect 258 -2 262 18
rect 266 -2 270 18
rect 404 19 408 59
rect 412 19 416 59
rect 426 19 430 59
rect 434 19 438 59
rect 449 19 453 59
rect 457 19 461 59
rect 471 19 475 59
rect 479 19 483 59
rect 503 42 508 62
rect 512 42 516 62
rect 542 42 547 62
rect 551 42 555 62
rect 568 40 572 60
rect 576 40 580 60
rect 584 40 588 60
rect 592 40 596 60
rect 298 7 318 11
rect 298 -1 318 3
rect 329 -9 333 11
rect 337 -9 341 11
rect 359 -2 363 18
rect 367 -2 371 18
rect -120 -47 -116 -27
rect -112 -47 -108 -27
rect -104 -47 -100 -27
rect -96 -47 -92 -27
rect 55 -34 75 -30
rect 55 -42 75 -38
rect 55 -59 75 -55
rect 55 -67 75 -63
rect 99 -72 103 -52
rect 107 -72 111 -52
rect 115 -72 119 -52
rect 123 -72 127 -52
rect 143 -72 147 -52
rect 151 -72 155 -52
rect 185 -70 189 -30
rect 193 -70 197 -30
rect 201 -70 205 -30
rect 209 -70 213 -30
rect 222 -70 226 -30
rect 230 -70 234 -30
rect 245 -70 249 -50
rect 253 -70 257 -50
rect 279 -70 283 -30
rect 287 -70 291 -30
rect 295 -70 299 -30
rect 303 -70 307 -30
rect 316 -70 320 -30
rect 324 -70 328 -30
rect 339 -70 343 -50
rect 347 -70 351 -50
rect 373 -70 377 -30
rect 381 -70 385 -30
rect 389 -70 393 -30
rect 397 -70 401 -30
rect 410 -70 414 -30
rect 418 -70 422 -30
rect 433 -70 437 -50
rect 441 -70 445 -50
rect -11 -106 -7 -86
rect -3 -106 1 -86
rect 19 -99 23 -79
rect 27 -99 31 -79
rect 42 -91 62 -87
rect 42 -99 62 -95
rect -284 -161 -280 -121
rect -276 -161 -272 -121
rect -262 -161 -258 -121
rect -254 -161 -250 -121
rect -239 -161 -235 -121
rect -231 -161 -227 -121
rect -217 -161 -213 -121
rect -209 -161 -205 -121
rect -185 -138 -180 -118
rect -176 -138 -172 -118
rect -146 -138 -141 -118
rect -137 -138 -133 -118
rect -120 -140 -116 -120
rect -112 -140 -108 -120
rect -104 -140 -100 -120
rect -96 -140 -92 -120
rect 457 -72 461 -32
rect 465 -72 469 -32
rect 479 -72 483 -32
rect 487 -72 491 -32
rect 502 -72 506 -32
rect 510 -72 514 -32
rect 524 -72 528 -32
rect 532 -72 536 -32
rect 556 -49 561 -29
rect 565 -49 569 -29
rect 595 -49 600 -29
rect 604 -49 608 -29
rect 621 -51 625 -31
rect 629 -51 633 -31
rect 637 -51 641 -31
rect 645 -51 649 -31
rect 36 -159 56 -155
rect 99 -160 103 -140
rect 107 -160 111 -140
rect 118 -160 122 -140
rect 126 -160 130 -140
rect 137 -160 141 -140
rect 145 -160 149 -140
rect 156 -160 160 -140
rect 164 -160 168 -140
rect 172 -160 176 -140
rect 180 -160 184 -140
rect 210 -156 214 -136
rect 218 -156 222 -136
rect 226 -156 230 -136
rect 234 -156 238 -136
rect 255 -156 259 -136
rect 263 -156 267 -136
rect 354 -155 374 -151
rect 36 -167 56 -163
rect 36 -175 56 -171
rect 354 -163 374 -159
rect 36 -183 56 -179
rect 36 -200 56 -196
rect 36 -208 56 -204
rect -284 -255 -280 -215
rect -276 -255 -272 -215
rect -262 -255 -258 -215
rect -254 -255 -250 -215
rect -239 -255 -235 -215
rect -231 -255 -227 -215
rect -217 -255 -213 -215
rect -209 -255 -205 -215
rect -185 -232 -180 -212
rect -176 -232 -172 -212
rect -146 -232 -141 -212
rect -137 -232 -133 -212
rect -120 -234 -116 -214
rect -112 -234 -108 -214
rect -104 -234 -100 -214
rect -96 -234 -92 -214
rect 354 -177 394 -173
rect 443 -177 447 -137
rect 451 -177 455 -137
rect 465 -177 469 -137
rect 473 -177 477 -137
rect 488 -177 492 -137
rect 496 -177 500 -137
rect 510 -177 514 -137
rect 518 -177 522 -137
rect 542 -180 547 -160
rect 551 -180 555 -160
rect 581 -180 586 -160
rect 590 -180 594 -160
rect 607 -178 611 -158
rect 615 -178 619 -158
rect 623 -178 627 -158
rect 631 -178 635 -158
rect 354 -185 394 -181
rect 354 -197 394 -193
rect 354 -205 394 -201
rect 453 -207 493 -203
rect 453 -215 493 -211
rect -28 -247 -24 -227
rect -20 -247 -16 -227
rect 2 -240 6 -220
rect 10 -240 14 -220
rect 25 -232 45 -228
rect 25 -240 45 -236
rect 107 -259 111 -239
rect 115 -259 119 -239
rect 126 -259 130 -239
rect 134 -259 138 -239
rect 145 -259 149 -239
rect 153 -259 157 -239
rect 164 -259 168 -239
rect 172 -259 176 -239
rect 180 -259 184 -239
rect 188 -259 192 -239
rect 210 -240 214 -220
rect 218 -240 222 -220
rect 226 -240 230 -220
rect 234 -240 238 -220
rect 249 -240 253 -220
rect 257 -240 261 -220
rect 274 -240 278 -220
rect 282 -240 286 -220
rect 453 -229 493 -225
rect 354 -233 374 -229
rect 453 -237 493 -233
rect 354 -241 374 -237
rect 354 -254 414 -250
rect 453 -252 493 -248
rect 19 -300 39 -296
rect -284 -349 -280 -309
rect -276 -349 -272 -309
rect -262 -349 -258 -309
rect -254 -349 -250 -309
rect -239 -349 -235 -309
rect -231 -349 -227 -309
rect -217 -349 -213 -309
rect -209 -349 -205 -309
rect -185 -326 -180 -306
rect -176 -326 -172 -306
rect -146 -326 -141 -306
rect -137 -326 -133 -306
rect 19 -308 39 -304
rect -120 -328 -116 -308
rect -112 -328 -108 -308
rect -104 -328 -100 -308
rect -96 -328 -92 -308
rect 19 -316 39 -312
rect 354 -262 414 -258
rect 453 -260 493 -256
rect 354 -275 414 -271
rect 453 -274 493 -270
rect 354 -283 414 -279
rect 453 -282 493 -278
rect 354 -296 414 -292
rect 354 -304 414 -300
rect 450 -307 470 -302
rect 19 -324 39 -320
rect 210 -334 214 -314
rect 218 -334 222 -314
rect 226 -334 230 -314
rect 234 -334 238 -314
rect 251 -334 255 -314
rect 259 -334 263 -314
rect 279 -334 283 -314
rect 287 -334 291 -314
rect 450 -315 470 -311
rect 19 -341 39 -337
rect 19 -349 39 -345
rect 111 -359 115 -339
rect 119 -359 123 -339
rect 127 -359 131 -339
rect 135 -359 139 -339
rect 150 -359 154 -339
rect 158 -359 162 -339
rect 175 -359 179 -339
rect 183 -359 187 -339
rect 356 -341 376 -337
rect 356 -349 376 -345
rect 450 -346 470 -341
rect -46 -388 -42 -368
rect -38 -388 -34 -368
rect -16 -381 -12 -361
rect -8 -381 -4 -361
rect 7 -373 27 -369
rect 7 -381 27 -377
rect -284 -443 -280 -403
rect -276 -443 -272 -403
rect -262 -443 -258 -403
rect -254 -443 -250 -403
rect -239 -443 -235 -403
rect -231 -443 -227 -403
rect -217 -443 -213 -403
rect -209 -443 -205 -403
rect -185 -420 -180 -400
rect -176 -420 -172 -400
rect -146 -420 -141 -400
rect -137 -420 -133 -400
rect -120 -422 -116 -402
rect -112 -422 -108 -402
rect -104 -422 -100 -402
rect -96 -422 -92 -402
rect 450 -354 470 -350
rect 356 -363 436 -359
rect 356 -371 436 -367
rect 452 -371 472 -367
rect 452 -379 472 -375
rect 356 -385 436 -381
rect 452 -387 472 -383
rect 356 -393 436 -389
rect 452 -395 472 -391
rect 356 -407 436 -403
rect 210 -428 214 -408
rect 218 -428 222 -408
rect 226 -428 230 -408
rect 234 -428 238 -408
rect 251 -428 255 -408
rect 259 -428 263 -408
rect 356 -415 436 -411
rect 1 -441 21 -437
rect 1 -449 21 -445
rect 104 -453 108 -433
rect 112 -453 116 -433
rect 120 -453 124 -433
rect 128 -453 132 -433
rect 145 -453 149 -433
rect 153 -453 157 -433
rect 356 -428 436 -424
rect 356 -436 436 -432
rect 1 -457 21 -453
rect 1 -465 21 -461
rect 1 -482 21 -478
rect 1 -490 21 -486
<< polysilicon >>
rect -179 163 -177 166
rect -140 163 -138 166
rect -279 160 -277 163
rect -257 160 -255 163
rect -234 160 -232 163
rect -212 160 -210 163
rect -115 161 -113 164
rect -99 161 -97 164
rect 44 163 46 166
rect 83 163 85 166
rect -179 141 -177 143
rect -140 141 -138 143
rect -56 160 -54 163
rect -34 160 -32 163
rect -11 160 -9 163
rect 11 160 13 163
rect -179 139 -169 141
rect -140 139 -130 141
rect -279 104 -277 120
rect -257 99 -255 120
rect -234 104 -232 120
rect -212 99 -210 120
rect -188 119 -186 128
rect -171 127 -169 139
rect -171 119 -169 122
rect -149 119 -147 128
rect -132 127 -130 139
rect -132 119 -130 122
rect -115 120 -113 141
rect -99 120 -97 141
rect 108 161 110 164
rect 124 161 126 164
rect 44 141 46 143
rect 83 141 85 143
rect 499 158 501 161
rect 538 158 540 161
rect 399 155 401 158
rect 421 155 423 158
rect 444 155 446 158
rect 466 155 468 158
rect 44 139 54 141
rect 83 139 93 141
rect -115 113 -113 116
rect -99 113 -97 116
rect -56 104 -54 120
rect -188 96 -186 99
rect -171 95 -169 99
rect -149 96 -147 99
rect -132 95 -130 99
rect -34 99 -32 120
rect -11 104 -9 120
rect 11 99 13 120
rect 35 119 37 128
rect 52 127 54 139
rect 52 119 54 122
rect 74 119 76 128
rect 91 127 93 139
rect 91 119 93 122
rect 108 120 110 141
rect 124 120 126 141
rect 262 116 264 119
rect 364 116 366 119
rect 108 113 110 116
rect 124 113 126 116
rect 232 108 234 111
rect 193 102 196 104
rect 206 102 213 104
rect 35 96 37 99
rect 52 95 54 99
rect 74 96 76 99
rect 91 95 93 99
rect -279 91 -277 94
rect -234 91 -232 94
rect -56 91 -54 94
rect -11 91 -9 94
rect 232 83 234 98
rect 262 90 264 106
rect 334 108 336 111
rect 295 102 298 104
rect 308 102 315 104
rect 563 156 565 159
rect 579 156 581 159
rect 499 136 501 138
rect 538 136 540 138
rect 499 134 509 136
rect 538 134 548 136
rect 193 76 196 78
rect 216 76 223 78
rect -179 69 -177 72
rect -140 69 -138 72
rect -279 66 -277 69
rect -257 66 -255 69
rect -234 66 -232 69
rect -212 66 -210 69
rect -115 67 -113 70
rect -99 67 -97 70
rect -179 47 -177 49
rect -140 47 -138 49
rect 43 62 45 65
rect 334 83 336 98
rect 364 90 366 106
rect 399 99 401 115
rect 295 76 298 78
rect 318 76 325 78
rect 262 67 264 70
rect 421 94 423 115
rect 444 99 446 115
rect 466 94 468 115
rect 490 114 492 123
rect 507 122 509 134
rect 507 114 509 117
rect 529 114 531 123
rect 546 122 548 134
rect 546 114 548 117
rect 563 115 565 136
rect 579 115 581 136
rect 563 108 565 111
rect 579 108 581 111
rect 490 91 492 94
rect 507 90 509 94
rect 529 91 531 94
rect 546 90 548 94
rect 399 86 401 89
rect 444 86 446 89
rect 364 67 366 70
rect 13 55 15 58
rect -179 45 -169 47
rect -140 45 -130 47
rect -279 10 -277 26
rect -257 5 -255 26
rect -234 10 -232 26
rect -212 5 -210 26
rect -188 25 -186 34
rect -171 33 -169 45
rect -171 25 -169 28
rect -149 25 -147 34
rect -132 33 -130 45
rect -132 25 -130 28
rect -115 26 -113 47
rect -99 26 -97 47
rect 232 60 234 63
rect 334 60 336 63
rect 509 62 511 65
rect 548 62 550 65
rect 409 59 411 62
rect 431 59 433 62
rect 454 59 456 62
rect 476 59 478 62
rect 106 49 108 52
rect 122 49 124 52
rect 143 49 145 52
rect 54 47 61 49
rect 81 47 84 49
rect -115 19 -113 22
rect -99 19 -97 22
rect 13 19 15 35
rect 43 27 45 42
rect 64 21 71 23
rect 81 21 84 23
rect 43 14 45 17
rect 263 44 265 47
rect 364 44 366 47
rect 233 36 235 39
rect 166 29 168 32
rect 194 30 197 32
rect 207 30 214 32
rect 233 11 235 26
rect 263 18 265 34
rect 334 36 336 39
rect 295 30 298 32
rect 308 30 315 32
rect 13 6 15 9
rect -188 2 -186 5
rect -171 1 -169 5
rect -149 2 -147 5
rect -132 1 -130 5
rect -279 -3 -277 0
rect -234 -3 -232 0
rect 106 -7 108 9
rect 122 -7 124 9
rect 16 -21 19 -19
rect 39 -21 55 -19
rect 75 -21 78 -19
rect -179 -25 -177 -22
rect -140 -25 -138 -22
rect -279 -28 -277 -25
rect -257 -28 -255 -25
rect -234 -28 -232 -25
rect -212 -28 -210 -25
rect -115 -27 -113 -24
rect -99 -27 -97 -24
rect 143 -21 145 9
rect 166 -7 168 9
rect 194 4 197 6
rect 217 4 224 6
rect 334 11 336 26
rect 364 18 366 34
rect 573 60 575 63
rect 589 60 591 63
rect 509 40 511 42
rect 548 40 550 42
rect 509 38 519 40
rect 548 38 558 40
rect 295 4 298 6
rect 318 4 325 6
rect 263 -5 265 -2
rect 409 3 411 19
rect 364 -5 366 -2
rect 431 -2 433 19
rect 454 3 456 19
rect 476 -2 478 19
rect 500 18 502 27
rect 517 26 519 38
rect 517 18 519 21
rect 539 18 541 27
rect 556 26 558 38
rect 556 18 558 21
rect 573 19 575 40
rect 589 19 591 40
rect 573 12 575 15
rect 589 12 591 15
rect 500 -5 502 -2
rect 517 -6 519 -2
rect 539 -5 541 -2
rect 556 -6 558 -2
rect 233 -12 235 -9
rect 334 -12 336 -9
rect 409 -10 411 -7
rect 454 -10 456 -7
rect 166 -20 168 -17
rect -179 -47 -177 -45
rect -140 -47 -138 -45
rect 106 -30 108 -27
rect 122 -30 124 -27
rect 190 -30 192 -27
rect 206 -30 208 -27
rect 227 -30 229 -27
rect 284 -30 286 -27
rect 300 -30 302 -27
rect 321 -30 323 -27
rect 378 -30 380 -27
rect 394 -30 396 -27
rect 415 -30 417 -27
rect 562 -29 564 -26
rect 601 -29 603 -26
rect 143 -35 145 -31
rect 16 -37 19 -35
rect 39 -37 55 -35
rect 75 -37 78 -35
rect -179 -49 -169 -47
rect -140 -49 -130 -47
rect -279 -84 -277 -68
rect -257 -89 -255 -68
rect -234 -84 -232 -68
rect -212 -89 -210 -68
rect -188 -69 -186 -60
rect -171 -61 -169 -49
rect -171 -69 -169 -66
rect -149 -69 -147 -60
rect -132 -61 -130 -49
rect -132 -69 -130 -66
rect -115 -68 -113 -47
rect -99 -68 -97 -47
rect 104 -52 106 -49
rect 120 -52 122 -49
rect 148 -52 150 -49
rect 26 -62 29 -60
rect 39 -62 55 -60
rect 75 -62 78 -60
rect 250 -50 252 -47
rect 344 -50 346 -47
rect 462 -32 464 -29
rect 484 -32 486 -29
rect 507 -32 509 -29
rect 529 -32 531 -29
rect 438 -50 440 -47
rect -115 -75 -113 -72
rect -99 -75 -97 -72
rect 24 -79 26 -76
rect -6 -86 -4 -83
rect -188 -92 -186 -89
rect -171 -93 -169 -89
rect -149 -92 -147 -89
rect -132 -93 -130 -89
rect -279 -97 -277 -94
rect -234 -97 -232 -94
rect 104 -88 106 -72
rect 120 -88 122 -72
rect 148 -88 150 -72
rect 190 -86 192 -70
rect 206 -86 208 -70
rect 35 -94 42 -92
rect 62 -94 65 -92
rect -179 -118 -177 -115
rect -140 -118 -138 -115
rect -279 -121 -277 -118
rect -257 -121 -255 -118
rect -234 -121 -232 -118
rect -212 -121 -210 -118
rect -115 -120 -113 -117
rect -99 -120 -97 -117
rect -179 -140 -177 -138
rect -140 -140 -138 -138
rect -6 -122 -4 -106
rect 24 -114 26 -99
rect 148 -101 150 -98
rect 227 -100 229 -70
rect 250 -86 252 -70
rect 284 -86 286 -70
rect 300 -86 302 -70
rect 250 -99 252 -96
rect 104 -111 106 -108
rect 120 -111 122 -108
rect 190 -109 192 -106
rect 206 -109 208 -106
rect 321 -100 323 -70
rect 344 -86 346 -70
rect 378 -86 380 -70
rect 394 -86 396 -70
rect 344 -99 346 -96
rect 284 -109 286 -106
rect 300 -109 302 -106
rect 415 -100 417 -70
rect 438 -86 440 -70
rect 626 -31 628 -28
rect 642 -31 644 -28
rect 562 -51 564 -49
rect 601 -51 603 -49
rect 562 -53 572 -51
rect 601 -53 611 -51
rect 462 -88 464 -72
rect 438 -99 440 -96
rect 484 -93 486 -72
rect 507 -88 509 -72
rect 529 -93 531 -72
rect 553 -73 555 -64
rect 570 -65 572 -53
rect 570 -73 572 -70
rect 592 -73 594 -64
rect 609 -65 611 -53
rect 609 -73 611 -70
rect 626 -72 628 -51
rect 642 -72 644 -51
rect 626 -79 628 -76
rect 642 -79 644 -76
rect 553 -96 555 -93
rect 570 -97 572 -93
rect 592 -96 594 -93
rect 609 -97 611 -93
rect 378 -109 380 -106
rect 394 -109 396 -106
rect 462 -101 464 -98
rect 507 -101 509 -98
rect 227 -114 229 -110
rect 321 -114 323 -110
rect 415 -114 417 -110
rect 448 -111 450 -108
rect 493 -111 495 -108
rect 45 -120 52 -118
rect 62 -120 65 -118
rect 24 -127 26 -124
rect -6 -135 -4 -132
rect 215 -136 217 -133
rect 231 -136 233 -133
rect 260 -136 262 -133
rect 104 -140 106 -137
rect 123 -140 125 -137
rect 142 -140 144 -137
rect 161 -140 163 -137
rect 177 -140 179 -137
rect -179 -142 -169 -140
rect -140 -142 -130 -140
rect -279 -177 -277 -161
rect -257 -182 -255 -161
rect -234 -177 -232 -161
rect -212 -182 -210 -161
rect -188 -162 -186 -153
rect -171 -154 -169 -142
rect -171 -162 -169 -159
rect -149 -162 -147 -153
rect -132 -154 -130 -142
rect -132 -162 -130 -159
rect -115 -161 -113 -140
rect -99 -161 -97 -140
rect 448 -137 450 -121
rect 470 -137 472 -116
rect 539 -116 541 -113
rect 556 -116 558 -112
rect 578 -116 580 -113
rect 595 -116 597 -112
rect 493 -137 495 -121
rect 515 -137 517 -116
rect 612 -133 614 -130
rect 628 -133 630 -130
rect -3 -162 0 -160
rect 20 -162 36 -160
rect 56 -162 59 -160
rect -115 -168 -113 -165
rect -99 -168 -97 -165
rect -3 -178 0 -176
rect 20 -178 36 -176
rect 56 -178 59 -176
rect 104 -177 106 -160
rect 123 -177 125 -160
rect 142 -177 144 -160
rect 161 -177 163 -160
rect 177 -174 179 -160
rect 215 -172 217 -156
rect 231 -172 233 -156
rect 260 -172 262 -156
rect 325 -158 328 -156
rect 338 -158 354 -156
rect 374 -158 377 -156
rect -188 -185 -186 -182
rect -171 -186 -169 -182
rect -149 -185 -147 -182
rect -132 -186 -130 -182
rect -279 -190 -277 -187
rect -234 -190 -232 -187
rect 7 -203 10 -201
rect 20 -203 36 -201
rect 56 -203 59 -201
rect -179 -212 -177 -209
rect -140 -212 -138 -209
rect -279 -215 -277 -212
rect -257 -215 -255 -212
rect -234 -215 -232 -212
rect -212 -215 -210 -212
rect -115 -214 -113 -211
rect -99 -214 -97 -211
rect -179 -234 -177 -232
rect -140 -234 -138 -232
rect 177 -187 179 -184
rect 539 -145 541 -136
rect 556 -139 558 -136
rect 556 -156 558 -144
rect 578 -145 580 -136
rect 595 -139 597 -136
rect 595 -156 597 -144
rect 548 -158 558 -156
rect 587 -158 597 -156
rect 612 -158 614 -137
rect 628 -158 630 -137
rect 548 -160 550 -158
rect 587 -160 589 -158
rect 325 -180 328 -178
rect 338 -180 354 -178
rect 394 -180 397 -178
rect 448 -180 450 -177
rect 470 -180 472 -177
rect 493 -180 495 -177
rect 515 -180 517 -177
rect 260 -185 262 -182
rect 548 -183 550 -180
rect 587 -183 589 -180
rect 612 -181 614 -178
rect 628 -181 630 -178
rect 215 -195 217 -192
rect 231 -195 233 -192
rect 325 -200 328 -198
rect 338 -200 354 -198
rect 394 -200 397 -198
rect 450 -210 453 -208
rect 493 -210 509 -208
rect 519 -210 522 -208
rect 7 -220 9 -217
rect -23 -227 -21 -224
rect -179 -236 -169 -234
rect -140 -236 -130 -234
rect -279 -271 -277 -255
rect -257 -276 -255 -255
rect -234 -271 -232 -255
rect -212 -276 -210 -255
rect -188 -256 -186 -247
rect -171 -248 -169 -236
rect -171 -256 -169 -253
rect -149 -256 -147 -247
rect -132 -248 -130 -236
rect -132 -256 -130 -253
rect -115 -255 -113 -234
rect -99 -255 -97 -234
rect 104 -221 106 -217
rect 123 -221 125 -217
rect 142 -221 144 -217
rect 161 -221 163 -217
rect 215 -220 217 -217
rect 231 -220 233 -217
rect 254 -220 256 -217
rect 279 -220 281 -217
rect 18 -235 25 -233
rect 45 -235 48 -233
rect 112 -239 114 -236
rect 131 -239 133 -236
rect 150 -239 152 -236
rect 169 -239 171 -236
rect 185 -239 187 -236
rect -115 -262 -113 -259
rect -99 -262 -97 -259
rect -23 -263 -21 -247
rect 7 -255 9 -240
rect 450 -232 453 -230
rect 493 -232 514 -230
rect 325 -236 328 -234
rect 338 -236 354 -234
rect 374 -236 377 -234
rect 215 -256 217 -240
rect 231 -256 233 -240
rect 254 -256 256 -240
rect 279 -256 281 -240
rect 450 -255 453 -253
rect 493 -255 509 -253
rect 519 -255 522 -253
rect 28 -261 35 -259
rect 45 -261 48 -259
rect 7 -268 9 -265
rect -23 -276 -21 -273
rect 112 -276 114 -259
rect 131 -276 133 -259
rect 150 -276 152 -259
rect 169 -276 171 -259
rect 185 -273 187 -259
rect -188 -279 -186 -276
rect -171 -280 -169 -276
rect -149 -279 -147 -276
rect -132 -280 -130 -276
rect -279 -284 -277 -281
rect -234 -284 -232 -281
rect -20 -303 -17 -301
rect 3 -303 19 -301
rect 39 -303 42 -301
rect -179 -306 -177 -303
rect -140 -306 -138 -303
rect -279 -309 -277 -306
rect -257 -309 -255 -306
rect -234 -309 -232 -306
rect -212 -309 -210 -306
rect -115 -308 -113 -305
rect -99 -308 -97 -305
rect -179 -328 -177 -326
rect -140 -328 -138 -326
rect 185 -286 187 -283
rect 325 -257 328 -255
rect 338 -257 354 -255
rect 414 -257 417 -255
rect 279 -269 281 -266
rect 325 -278 328 -276
rect 338 -278 354 -276
rect 414 -278 417 -276
rect 450 -277 453 -275
rect 493 -277 514 -275
rect 215 -289 217 -286
rect 231 -289 233 -286
rect 254 -289 256 -286
rect 325 -299 328 -297
rect 338 -299 354 -297
rect 414 -299 417 -297
rect 485 -301 494 -299
rect 514 -301 517 -299
rect 447 -310 450 -308
rect 470 -310 474 -308
rect 215 -314 217 -311
rect 231 -314 233 -311
rect 256 -314 258 -311
rect 284 -314 286 -311
rect -20 -319 -17 -317
rect 3 -319 19 -317
rect 39 -319 42 -317
rect 112 -320 114 -316
rect 131 -320 133 -316
rect 150 -320 152 -316
rect 169 -320 171 -316
rect -179 -330 -169 -328
rect -140 -330 -130 -328
rect -279 -365 -277 -349
rect -257 -370 -255 -349
rect -234 -365 -232 -349
rect -212 -370 -210 -349
rect -188 -350 -186 -341
rect -171 -342 -169 -330
rect -171 -350 -169 -347
rect -149 -350 -147 -341
rect -132 -342 -130 -330
rect -132 -350 -130 -347
rect -115 -349 -113 -328
rect -99 -349 -97 -328
rect 472 -316 474 -310
rect 472 -318 486 -316
rect 491 -318 494 -316
rect 514 -318 518 -316
rect 116 -339 118 -336
rect 132 -339 134 -336
rect 155 -339 157 -336
rect 180 -339 182 -336
rect -10 -344 -7 -342
rect 3 -344 19 -342
rect 39 -344 42 -342
rect -115 -356 -113 -353
rect -99 -356 -97 -353
rect -11 -361 -9 -358
rect 215 -350 217 -334
rect 231 -350 233 -334
rect 256 -350 258 -334
rect 284 -350 286 -334
rect 485 -340 494 -338
rect 514 -340 517 -338
rect 327 -344 330 -342
rect 340 -344 356 -342
rect 376 -344 379 -342
rect 447 -349 450 -347
rect 470 -349 474 -347
rect -41 -368 -39 -365
rect -188 -373 -186 -370
rect -171 -374 -169 -370
rect -149 -373 -147 -370
rect -132 -374 -130 -370
rect -279 -378 -277 -375
rect -234 -378 -232 -375
rect 0 -376 7 -374
rect 27 -376 30 -374
rect 116 -375 118 -359
rect 132 -375 134 -359
rect 155 -375 157 -359
rect 180 -375 182 -359
rect -179 -400 -177 -397
rect -140 -400 -138 -397
rect -279 -403 -277 -400
rect -257 -403 -255 -400
rect -234 -403 -232 -400
rect -212 -403 -210 -400
rect -115 -402 -113 -399
rect -99 -402 -97 -399
rect -179 -422 -177 -420
rect -140 -422 -138 -420
rect -41 -404 -39 -388
rect -11 -396 -9 -381
rect 10 -402 17 -400
rect 27 -402 30 -400
rect -11 -409 -9 -406
rect 472 -355 474 -349
rect 472 -357 486 -355
rect 284 -363 286 -360
rect 491 -357 494 -355
rect 514 -357 518 -355
rect 327 -366 330 -364
rect 340 -366 356 -364
rect 436 -366 439 -364
rect 449 -374 452 -372
rect 472 -374 493 -372
rect 497 -374 500 -372
rect 215 -383 217 -380
rect 231 -383 233 -380
rect 256 -383 258 -380
rect 180 -388 182 -385
rect 327 -388 330 -386
rect 340 -388 356 -386
rect 436 -388 439 -386
rect 449 -390 452 -388
rect 472 -390 493 -388
rect 497 -390 500 -388
rect 116 -408 118 -405
rect 132 -408 134 -405
rect 155 -408 157 -405
rect 215 -408 217 -405
rect 231 -408 233 -405
rect 256 -408 258 -405
rect -41 -417 -39 -414
rect -179 -424 -169 -422
rect -140 -424 -130 -422
rect -279 -459 -277 -443
rect -257 -464 -255 -443
rect -234 -459 -232 -443
rect -212 -464 -210 -443
rect -188 -444 -186 -435
rect -171 -436 -169 -424
rect -171 -444 -169 -441
rect -149 -444 -147 -435
rect -132 -436 -130 -424
rect -132 -444 -130 -441
rect -115 -443 -113 -422
rect -99 -443 -97 -422
rect 327 -410 330 -408
rect 340 -410 356 -408
rect 436 -410 439 -408
rect 109 -433 111 -430
rect 125 -433 127 -430
rect 150 -433 152 -430
rect -38 -444 -35 -442
rect -15 -444 1 -442
rect 21 -444 24 -442
rect -115 -450 -113 -447
rect -99 -450 -97 -447
rect 215 -444 217 -428
rect 231 -444 233 -428
rect 256 -444 258 -428
rect 327 -431 330 -429
rect 340 -431 356 -429
rect 436 -431 439 -429
rect -38 -460 -35 -458
rect -15 -460 1 -458
rect 21 -460 24 -458
rect -188 -467 -186 -464
rect -171 -468 -169 -464
rect -149 -467 -147 -464
rect -132 -468 -130 -464
rect 109 -469 111 -453
rect 125 -469 127 -453
rect 150 -469 152 -453
rect 256 -457 258 -454
rect 215 -467 217 -464
rect 231 -467 233 -464
rect -279 -472 -277 -469
rect -234 -472 -232 -469
rect -28 -485 -25 -483
rect -15 -485 1 -483
rect 21 -485 24 -483
rect 150 -482 152 -479
rect 109 -492 111 -489
rect 125 -492 127 -489
<< polycontact >>
rect -193 122 -188 127
rect -283 107 -279 111
rect -261 99 -257 104
rect -238 107 -234 111
rect -216 99 -212 104
rect -171 122 -167 127
rect -153 122 -149 127
rect -119 129 -115 133
rect -132 122 -128 127
rect -103 129 -99 133
rect 30 122 35 127
rect -60 107 -56 111
rect -38 99 -34 104
rect -15 107 -11 111
rect 7 99 11 104
rect 52 122 56 127
rect 70 122 74 127
rect 104 129 108 133
rect 91 122 95 127
rect 120 129 124 133
rect 209 104 213 108
rect 234 91 238 95
rect 311 104 315 108
rect 264 98 268 102
rect 485 117 490 122
rect 219 72 223 76
rect 336 91 340 95
rect 395 102 399 106
rect 366 98 370 102
rect 321 72 325 76
rect 417 94 421 99
rect 440 102 444 106
rect 462 94 466 99
rect 507 117 511 122
rect 525 117 529 122
rect 559 124 563 128
rect 546 117 550 122
rect 575 124 579 128
rect -193 28 -188 33
rect -283 13 -279 17
rect -261 5 -257 10
rect -238 13 -234 17
rect -216 5 -212 10
rect -171 28 -167 33
rect -153 28 -149 33
rect -119 35 -115 39
rect -132 28 -128 33
rect -103 35 -99 39
rect 54 49 58 53
rect 9 23 13 27
rect 39 30 43 34
rect 64 17 68 21
rect 210 32 214 36
rect 235 19 239 23
rect 311 32 315 36
rect 265 26 269 30
rect 102 -4 106 0
rect 124 -4 128 0
rect 42 -19 46 -15
rect 162 -4 166 0
rect 220 0 224 4
rect 145 -18 149 -14
rect 336 19 340 23
rect 366 26 370 30
rect 495 21 500 26
rect 321 0 325 4
rect 405 6 409 10
rect 427 -2 431 3
rect 450 6 454 10
rect 472 -2 476 3
rect 517 21 521 26
rect 535 21 539 26
rect 569 28 573 32
rect 556 21 560 26
rect 585 28 589 32
rect 42 -41 46 -37
rect -193 -66 -188 -61
rect -283 -81 -279 -77
rect -261 -89 -257 -84
rect -238 -81 -234 -77
rect -216 -89 -212 -84
rect -171 -66 -167 -61
rect -153 -66 -149 -61
rect -119 -59 -115 -55
rect -132 -66 -128 -61
rect -103 -59 -99 -55
rect 42 -60 46 -56
rect 100 -85 104 -81
rect 35 -92 39 -88
rect 122 -85 126 -81
rect 144 -85 148 -81
rect 186 -83 190 -79
rect 208 -83 212 -79
rect -10 -118 -6 -114
rect 20 -111 24 -107
rect 246 -83 250 -79
rect 280 -83 284 -79
rect 302 -83 306 -79
rect 229 -97 233 -93
rect 340 -83 344 -79
rect 374 -83 378 -79
rect 396 -83 400 -79
rect 323 -97 327 -93
rect 434 -83 438 -79
rect 548 -70 553 -65
rect 458 -85 462 -81
rect 417 -97 421 -93
rect 480 -93 484 -88
rect 503 -85 507 -81
rect 525 -93 529 -88
rect 570 -70 574 -65
rect 588 -70 592 -65
rect 622 -63 626 -59
rect 609 -70 613 -65
rect 638 -63 642 -59
rect 45 -124 49 -120
rect 466 -121 470 -116
rect 444 -128 448 -124
rect -193 -159 -188 -154
rect -283 -174 -279 -170
rect -261 -182 -257 -177
rect -238 -174 -234 -170
rect -216 -182 -212 -177
rect -171 -159 -167 -154
rect -153 -159 -149 -154
rect -119 -152 -115 -148
rect -132 -159 -128 -154
rect -103 -152 -99 -148
rect 23 -160 27 -156
rect 511 -121 515 -116
rect 489 -128 493 -124
rect 100 -173 104 -169
rect 119 -173 123 -169
rect 138 -173 142 -169
rect 157 -173 161 -169
rect 173 -171 177 -167
rect 211 -169 215 -165
rect 233 -169 237 -165
rect 256 -169 260 -165
rect 341 -163 346 -158
rect 23 -182 27 -178
rect 23 -201 27 -197
rect 534 -144 539 -139
rect 556 -144 560 -139
rect 574 -144 578 -139
rect 595 -144 599 -139
rect 608 -150 612 -146
rect 624 -150 628 -146
rect 341 -184 345 -180
rect 341 -204 345 -200
rect 502 -208 506 -204
rect -193 -253 -188 -248
rect -283 -268 -279 -264
rect -261 -276 -257 -271
rect -238 -268 -234 -264
rect -216 -276 -212 -271
rect -171 -253 -167 -248
rect -153 -253 -149 -248
rect -119 -246 -115 -242
rect -132 -253 -128 -248
rect -103 -246 -99 -242
rect 18 -233 22 -229
rect -27 -259 -23 -255
rect 3 -252 7 -248
rect 509 -230 514 -226
rect 211 -253 215 -249
rect 233 -253 237 -249
rect 256 -253 260 -249
rect 275 -253 279 -249
rect 341 -241 346 -236
rect 502 -253 506 -249
rect 28 -265 32 -261
rect 108 -272 112 -268
rect 127 -272 131 -268
rect 146 -272 150 -268
rect 165 -272 169 -268
rect 181 -270 185 -266
rect 6 -301 10 -297
rect 341 -261 345 -257
rect 509 -275 514 -271
rect 341 -282 345 -278
rect 486 -299 491 -294
rect 341 -303 345 -299
rect 6 -323 10 -319
rect -193 -347 -188 -342
rect -283 -362 -279 -358
rect -261 -370 -257 -365
rect -238 -362 -234 -358
rect -216 -370 -212 -365
rect -171 -347 -167 -342
rect -153 -347 -149 -342
rect -119 -340 -115 -336
rect -132 -347 -128 -342
rect -103 -340 -99 -336
rect 486 -320 491 -316
rect 6 -342 10 -338
rect 211 -347 215 -343
rect 233 -347 237 -343
rect 258 -347 262 -343
rect 280 -347 284 -343
rect 486 -338 491 -334
rect 343 -349 348 -344
rect 0 -374 4 -370
rect 112 -372 116 -368
rect 134 -372 138 -368
rect 157 -372 161 -368
rect 176 -372 180 -368
rect -45 -400 -41 -396
rect -15 -393 -11 -389
rect 10 -406 14 -402
rect 486 -359 491 -355
rect 343 -370 347 -366
rect 480 -372 484 -368
rect 480 -388 484 -384
rect 343 -392 347 -388
rect -193 -441 -188 -436
rect -283 -456 -279 -452
rect -261 -464 -257 -459
rect -238 -456 -234 -452
rect -216 -464 -212 -459
rect -171 -441 -167 -436
rect -153 -441 -149 -436
rect -119 -434 -115 -430
rect -132 -441 -128 -436
rect -103 -434 -99 -430
rect 343 -414 347 -410
rect -12 -442 -8 -438
rect 211 -441 215 -437
rect 233 -441 237 -437
rect 252 -441 256 -437
rect 343 -435 347 -431
rect -12 -464 -8 -460
rect 105 -466 109 -462
rect 127 -466 131 -462
rect 146 -466 150 -462
rect -12 -483 -8 -479
<< metal1 >>
rect -290 169 135 173
rect -284 160 -280 169
rect -239 160 -235 169
rect -176 163 -171 169
rect -137 163 -132 169
rect -272 120 -271 160
rect -263 120 -262 160
rect -276 115 -258 120
rect -227 120 -226 160
rect -218 120 -217 160
rect -254 111 -250 120
rect -231 115 -213 120
rect -172 143 -171 163
rect -133 143 -132 163
rect -120 161 -116 169
rect -104 161 -100 169
rect -185 134 -180 143
rect -185 130 -167 134
rect -146 133 -141 143
rect -112 133 -108 141
rect -96 133 -92 141
rect -61 160 -57 169
rect -16 160 -12 169
rect 47 163 52 169
rect 86 163 91 169
rect -146 130 -119 133
rect -209 113 -205 120
rect -185 119 -180 130
rect -146 119 -141 130
rect -112 130 -103 133
rect -112 120 -108 130
rect -96 129 -88 133
rect -96 120 -92 129
rect -49 120 -48 160
rect -40 120 -39 160
rect -290 107 -283 111
rect -254 107 -238 111
rect -284 90 -280 94
rect -254 96 -250 107
rect -271 94 -250 96
rect -276 93 -250 94
rect -239 90 -235 94
rect -209 96 -205 108
rect -226 94 -205 96
rect -231 93 -205 94
rect -193 96 -189 99
rect -176 96 -172 99
rect -193 93 -172 96
rect -168 90 -163 99
rect -154 96 -150 99
rect -137 96 -133 99
rect -154 93 -133 96
rect -129 90 -124 99
rect -120 90 -116 116
rect -104 90 -100 116
rect -53 115 -35 120
rect -4 120 -3 160
rect 5 120 6 160
rect -31 111 -27 120
rect -8 115 10 120
rect 51 143 52 163
rect 90 143 91 163
rect 103 161 107 169
rect 119 161 123 169
rect 165 164 602 168
rect 38 134 43 143
rect 38 130 56 134
rect 77 133 82 143
rect 394 155 398 164
rect 439 155 443 164
rect 502 158 507 164
rect 541 158 546 164
rect 111 133 115 141
rect 127 133 131 141
rect 77 130 104 133
rect 14 113 18 120
rect 38 119 43 130
rect 77 119 82 130
rect 111 130 120 133
rect 111 120 115 130
rect 127 129 135 133
rect 127 120 131 129
rect 181 131 278 134
rect -67 107 -60 111
rect -31 107 -15 111
rect -61 90 -57 94
rect -31 96 -27 107
rect -48 94 -27 96
rect -53 93 -27 94
rect -16 90 -12 94
rect 14 96 18 108
rect -3 94 18 96
rect -8 93 18 94
rect 30 96 34 99
rect 47 96 51 99
rect 30 93 51 96
rect 55 90 60 99
rect 69 96 73 99
rect 86 96 90 99
rect 69 93 90 96
rect 94 90 99 99
rect 103 90 107 116
rect 119 90 123 116
rect -290 88 123 90
rect 181 88 184 131
rect 254 121 255 128
rect 274 125 278 131
rect 272 124 383 125
rect 265 121 383 124
rect 265 116 269 121
rect 274 120 281 121
rect 209 112 257 116
rect 188 105 196 109
rect 209 108 213 112
rect 235 108 239 112
rect 188 96 192 105
rect 206 97 223 101
rect -290 85 184 88
rect -290 75 -91 79
rect -284 66 -280 75
rect -239 66 -235 75
rect -176 69 -171 75
rect -137 69 -132 75
rect -272 26 -271 66
rect -263 26 -262 66
rect -276 21 -258 26
rect -227 26 -226 66
rect -218 26 -217 66
rect -254 17 -250 26
rect -231 21 -213 26
rect -172 49 -171 69
rect -133 49 -132 69
rect -120 67 -116 75
rect -104 67 -100 75
rect -185 40 -180 49
rect -185 36 -167 40
rect -146 39 -141 49
rect -112 39 -108 47
rect -96 39 -92 47
rect -146 36 -119 39
rect -209 19 -205 26
rect -185 25 -180 36
rect -146 25 -141 36
rect -112 36 -103 39
rect -112 26 -108 36
rect -96 35 -89 39
rect -96 26 -92 35
rect -290 13 -283 17
rect -254 13 -238 17
rect -284 -4 -280 0
rect -254 2 -250 13
rect -271 0 -250 2
rect -276 -1 -250 0
rect -239 -4 -235 0
rect -209 2 -205 14
rect -226 0 -205 2
rect -231 -1 -205 0
rect -193 2 -189 5
rect -176 2 -172 5
rect -193 -1 -172 2
rect -168 -4 -163 5
rect -154 2 -150 5
rect -137 2 -133 5
rect -154 -1 -133 2
rect -129 -4 -124 5
rect -120 -4 -116 22
rect -104 -4 -100 22
rect -290 -5 -86 -4
rect -69 -5 -65 85
rect 188 75 192 91
rect 220 95 223 97
rect 227 95 231 98
rect 220 91 231 95
rect 238 91 242 95
rect 220 83 223 91
rect 216 79 223 83
rect 227 83 231 91
rect 257 90 261 106
rect 188 71 196 75
rect 219 67 223 72
rect 26 62 42 63
rect 26 58 38 62
rect -2 36 8 41
rect 182 62 219 65
rect 239 63 251 67
rect 235 62 251 63
rect 265 63 269 70
rect 54 53 58 58
rect 81 50 89 54
rect 95 53 112 57
rect 117 53 179 57
rect -12 23 4 27
rect -290 -9 -65 -5
rect -290 -19 -92 -15
rect -284 -28 -280 -19
rect -239 -28 -235 -19
rect -176 -25 -171 -19
rect -137 -25 -132 -19
rect -272 -68 -271 -28
rect -263 -68 -262 -28
rect -276 -73 -258 -68
rect -227 -68 -226 -28
rect -218 -68 -217 -28
rect -254 -77 -250 -68
rect -231 -73 -213 -68
rect -172 -45 -171 -25
rect -133 -45 -132 -25
rect -120 -27 -116 -19
rect -104 -27 -100 -19
rect -185 -54 -180 -45
rect -185 -58 -167 -54
rect -146 -55 -141 -45
rect -112 -55 -108 -47
rect -96 -55 -92 -47
rect -69 -55 -65 -9
rect -4 -45 -1 23
rect 16 19 20 35
rect 46 34 50 42
rect 54 42 61 46
rect 54 34 57 42
rect 35 30 39 34
rect 46 30 57 34
rect 46 27 50 30
rect 54 28 57 30
rect 85 34 89 50
rect 101 49 105 53
rect 125 49 129 53
rect 54 24 71 28
rect 38 13 42 17
rect 20 9 41 13
rect 2 5 12 9
rect 54 8 58 24
rect 85 20 89 29
rect 64 13 68 17
rect 81 16 89 20
rect 55 5 58 8
rect 109 5 113 9
rect 117 5 121 9
rect 138 5 142 9
rect 2 -30 7 5
rect 55 2 90 5
rect 26 -1 52 2
rect 87 0 90 2
rect 109 4 121 5
rect 109 0 115 4
rect 49 -4 83 -1
rect 38 -9 46 -6
rect 15 -18 19 -14
rect 42 -15 46 -9
rect 79 -14 83 -4
rect 75 -18 83 -14
rect 39 -26 55 -22
rect 42 -29 46 -26
rect 2 -34 19 -30
rect 47 -34 55 -30
rect 2 -55 7 -34
rect 15 -42 19 -38
rect 79 -38 83 -18
rect 42 -45 46 -41
rect 75 -42 83 -38
rect 33 -48 46 -45
rect -146 -58 -119 -55
rect -209 -75 -205 -68
rect -185 -69 -180 -58
rect -146 -69 -141 -58
rect -112 -58 -103 -55
rect -112 -68 -108 -58
rect -96 -59 -88 -55
rect -96 -68 -92 -59
rect -69 -59 29 -55
rect 79 -55 83 -42
rect -290 -81 -283 -77
rect -254 -81 -238 -77
rect -284 -98 -280 -94
rect -254 -92 -250 -81
rect -271 -94 -250 -92
rect -276 -95 -250 -94
rect -239 -98 -235 -94
rect -209 -92 -205 -80
rect -226 -94 -205 -92
rect -231 -95 -205 -94
rect -193 -92 -189 -89
rect -176 -92 -172 -89
rect -193 -95 -172 -92
rect -168 -98 -163 -89
rect -154 -92 -150 -89
rect -137 -92 -133 -89
rect -154 -95 -133 -92
rect -129 -98 -124 -89
rect -120 -98 -116 -72
rect -104 -98 -100 -72
rect -290 -99 -86 -98
rect -69 -99 -65 -59
rect 75 -59 83 -55
rect 87 -4 102 0
rect 120 0 121 4
rect 161 29 165 53
rect 146 0 150 9
rect 169 0 173 9
rect 182 0 185 62
rect 266 59 269 63
rect 266 58 275 59
rect 265 55 275 58
rect 278 52 281 120
rect 367 116 371 121
rect 311 112 359 116
rect 290 105 298 109
rect 311 108 315 112
rect 337 108 341 112
rect 290 96 294 105
rect 308 97 325 101
rect 290 75 294 91
rect 322 95 325 97
rect 329 95 333 98
rect 322 91 333 95
rect 340 91 344 95
rect 322 83 325 91
rect 318 79 325 83
rect 329 83 333 91
rect 359 90 363 106
rect 290 71 298 75
rect 321 67 325 72
rect 341 63 353 67
rect 337 62 353 63
rect 367 62 371 70
rect 369 57 371 62
rect 380 85 383 121
rect 406 115 407 155
rect 415 115 416 155
rect 402 110 420 115
rect 451 115 452 155
rect 460 115 461 155
rect 424 106 428 115
rect 447 110 465 115
rect 506 138 507 158
rect 545 138 546 158
rect 558 156 562 164
rect 574 156 578 164
rect 493 129 498 138
rect 493 125 511 129
rect 532 128 537 138
rect 566 128 570 136
rect 582 128 586 136
rect 532 125 559 128
rect 469 108 473 115
rect 493 114 498 125
rect 532 114 537 125
rect 566 125 575 128
rect 566 115 570 125
rect 582 124 592 128
rect 582 115 586 124
rect 393 104 395 106
rect 388 102 395 104
rect 424 102 440 106
rect 394 85 398 89
rect 424 91 428 102
rect 407 89 428 91
rect 402 88 428 89
rect 439 85 443 89
rect 469 91 473 103
rect 452 89 473 91
rect 447 88 473 89
rect 485 91 489 94
rect 502 91 506 94
rect 485 88 506 91
rect 510 85 515 94
rect 524 91 528 94
rect 541 91 545 94
rect 524 88 545 91
rect 549 85 554 94
rect 558 85 562 111
rect 574 85 578 111
rect 380 80 592 85
rect 380 52 383 80
rect 597 72 602 164
rect 398 68 602 72
rect 267 49 281 52
rect 363 49 383 52
rect 266 44 270 49
rect 367 44 371 49
rect 210 40 258 44
rect 189 33 197 37
rect 210 36 214 40
rect 236 36 240 40
rect 189 24 193 33
rect 207 25 224 29
rect 128 -4 130 0
rect 146 -4 162 0
rect 169 -4 185 0
rect 189 3 193 19
rect 221 23 224 25
rect 311 40 359 44
rect 228 23 232 26
rect 221 19 232 23
rect 239 19 243 23
rect 221 11 224 19
rect 217 7 224 11
rect 228 11 232 19
rect 258 18 262 34
rect 290 33 298 37
rect 311 36 315 40
rect 337 36 341 40
rect 290 24 294 33
rect 308 25 325 29
rect 189 -1 197 3
rect 87 -7 90 -4
rect 146 -7 150 -4
rect 169 -7 173 -4
rect 39 -67 55 -63
rect 42 -71 46 -67
rect 42 -75 76 -71
rect 7 -79 23 -78
rect 7 -83 19 -79
rect -290 -103 -65 -99
rect -290 -112 -91 -108
rect -284 -121 -280 -112
rect -239 -121 -235 -112
rect -176 -118 -171 -112
rect -137 -118 -132 -112
rect -272 -161 -271 -121
rect -263 -161 -262 -121
rect -276 -166 -258 -161
rect -227 -161 -226 -121
rect -218 -161 -217 -121
rect -254 -170 -250 -161
rect -231 -166 -213 -161
rect -172 -138 -171 -118
rect -133 -138 -132 -118
rect -120 -120 -116 -112
rect -104 -120 -100 -112
rect -185 -147 -180 -138
rect -185 -151 -167 -147
rect -146 -148 -141 -138
rect -112 -148 -108 -140
rect -146 -151 -119 -148
rect -209 -168 -205 -161
rect -185 -162 -180 -151
rect -146 -162 -141 -151
rect -112 -151 -103 -148
rect -112 -161 -108 -151
rect -96 -161 -92 -140
rect -290 -174 -283 -170
rect -254 -174 -238 -170
rect -284 -191 -280 -187
rect -254 -185 -250 -174
rect -271 -187 -250 -185
rect -276 -188 -250 -187
rect -239 -191 -235 -187
rect -209 -185 -205 -173
rect -226 -187 -205 -185
rect -231 -188 -205 -187
rect -193 -185 -189 -182
rect -176 -185 -172 -182
rect -193 -188 -172 -185
rect -168 -191 -163 -182
rect -154 -185 -150 -182
rect -137 -185 -133 -182
rect -154 -188 -133 -185
rect -129 -191 -124 -182
rect -120 -191 -116 -165
rect -104 -191 -100 -165
rect -290 -192 -86 -191
rect -69 -192 -65 -103
rect -21 -105 -11 -100
rect 35 -88 39 -83
rect 62 -91 70 -87
rect -31 -118 -15 -114
rect -23 -186 -20 -118
rect -3 -122 1 -106
rect 27 -107 31 -99
rect 35 -99 42 -95
rect 35 -107 38 -99
rect 16 -111 20 -107
rect 27 -111 38 -107
rect 27 -114 31 -111
rect 35 -113 38 -111
rect 66 -107 70 -91
rect 35 -117 52 -113
rect 19 -128 23 -124
rect 1 -132 22 -128
rect -17 -136 -7 -132
rect 35 -133 39 -117
rect 66 -121 70 -112
rect 45 -128 49 -124
rect 62 -125 70 -121
rect 36 -136 39 -133
rect -17 -171 -12 -136
rect 36 -139 66 -136
rect 7 -142 33 -139
rect 30 -145 64 -142
rect 19 -150 27 -147
rect -4 -159 0 -155
rect 23 -156 27 -150
rect 60 -155 64 -145
rect 56 -159 64 -155
rect 20 -167 36 -163
rect 23 -170 27 -167
rect -17 -175 0 -171
rect 28 -175 36 -171
rect -290 -196 -65 -192
rect -17 -196 -12 -175
rect -4 -183 0 -179
rect 60 -179 64 -159
rect 23 -186 27 -182
rect 56 -183 64 -179
rect 14 -189 27 -186
rect -69 -200 10 -196
rect 60 -196 64 -183
rect -290 -206 -91 -202
rect -284 -215 -280 -206
rect -239 -215 -235 -206
rect -176 -212 -171 -206
rect -137 -212 -132 -206
rect -272 -255 -271 -215
rect -263 -255 -262 -215
rect -276 -260 -258 -255
rect -227 -255 -226 -215
rect -218 -255 -217 -215
rect -254 -264 -250 -255
rect -231 -260 -213 -255
rect -172 -232 -171 -212
rect -133 -232 -132 -212
rect -120 -214 -116 -206
rect -104 -214 -100 -206
rect -185 -241 -180 -232
rect -185 -245 -167 -241
rect -146 -242 -141 -232
rect -112 -242 -108 -234
rect -146 -245 -119 -242
rect -209 -262 -205 -255
rect -185 -256 -180 -245
rect -146 -256 -141 -245
rect -112 -245 -103 -242
rect -112 -255 -108 -245
rect -96 -255 -92 -234
rect -290 -268 -283 -264
rect -254 -268 -238 -264
rect -284 -285 -280 -281
rect -254 -279 -250 -268
rect -271 -281 -250 -279
rect -276 -282 -250 -281
rect -239 -285 -235 -281
rect -209 -279 -205 -267
rect -226 -281 -205 -279
rect -231 -282 -205 -281
rect -193 -279 -189 -276
rect -176 -279 -172 -276
rect -193 -282 -172 -279
rect -168 -285 -163 -276
rect -154 -279 -150 -276
rect -137 -279 -133 -276
rect -154 -282 -133 -279
rect -129 -285 -124 -276
rect -120 -285 -116 -259
rect -104 -285 -100 -259
rect -290 -287 -86 -285
rect -69 -287 -65 -200
rect 56 -200 64 -196
rect 20 -208 36 -204
rect 23 -212 27 -208
rect 23 -216 62 -212
rect -10 -220 6 -219
rect -10 -224 2 -220
rect -53 -255 -49 -236
rect -38 -246 -28 -241
rect 18 -229 22 -224
rect 58 -220 62 -216
rect 45 -232 53 -228
rect -53 -259 -32 -255
rect -290 -290 -65 -287
rect -290 -300 -88 -296
rect -284 -309 -280 -300
rect -239 -309 -235 -300
rect -176 -306 -171 -300
rect -137 -306 -132 -300
rect -272 -349 -271 -309
rect -263 -349 -262 -309
rect -276 -354 -258 -349
rect -227 -349 -226 -309
rect -218 -349 -217 -309
rect -254 -358 -250 -349
rect -231 -354 -213 -349
rect -172 -326 -171 -306
rect -133 -326 -132 -306
rect -120 -308 -116 -300
rect -104 -308 -100 -300
rect -185 -335 -180 -326
rect -185 -339 -167 -335
rect -146 -336 -141 -326
rect -112 -336 -108 -328
rect -96 -336 -92 -328
rect -69 -335 -65 -290
rect -40 -327 -37 -259
rect -20 -263 -16 -247
rect 10 -248 14 -240
rect 18 -240 25 -236
rect 18 -248 21 -240
rect -1 -252 3 -248
rect 10 -252 21 -248
rect 10 -255 14 -252
rect 18 -254 21 -252
rect 49 -248 53 -232
rect 18 -258 35 -254
rect 2 -269 6 -265
rect -16 -273 5 -269
rect -34 -277 -24 -273
rect 18 -274 22 -258
rect 49 -262 53 -253
rect 28 -269 32 -265
rect 45 -266 53 -262
rect 19 -277 22 -274
rect -34 -312 -29 -277
rect 19 -280 49 -277
rect -10 -283 16 -280
rect 13 -286 47 -283
rect 51 -284 54 -280
rect 2 -291 10 -288
rect -21 -300 -17 -296
rect 6 -297 10 -291
rect 43 -296 47 -286
rect 39 -300 47 -296
rect 3 -308 19 -304
rect 6 -311 10 -308
rect -34 -316 -17 -312
rect 11 -316 19 -312
rect -146 -339 -119 -336
rect -209 -356 -205 -349
rect -185 -350 -180 -339
rect -146 -350 -141 -339
rect -112 -339 -103 -336
rect -112 -349 -108 -339
rect -96 -340 -89 -336
rect -96 -349 -92 -340
rect -73 -337 -65 -335
rect -34 -337 -29 -316
rect -21 -324 -17 -320
rect 43 -320 47 -300
rect 6 -327 10 -323
rect 39 -324 47 -320
rect -3 -330 10 -327
rect -73 -340 -7 -337
rect -74 -341 -7 -340
rect 43 -337 47 -324
rect -290 -362 -283 -358
rect -254 -362 -238 -358
rect -284 -379 -280 -375
rect -254 -373 -250 -362
rect -271 -375 -250 -373
rect -276 -376 -250 -375
rect -239 -379 -235 -375
rect -209 -373 -205 -361
rect -226 -375 -205 -373
rect -231 -376 -205 -375
rect -193 -373 -189 -370
rect -176 -373 -172 -370
rect -193 -376 -172 -373
rect -168 -379 -163 -370
rect -154 -373 -150 -370
rect -137 -373 -133 -370
rect -154 -376 -133 -373
rect -129 -379 -124 -370
rect -74 -345 -65 -341
rect 39 -341 47 -337
rect -120 -379 -116 -353
rect -104 -379 -100 -353
rect -290 -381 -86 -379
rect -74 -381 -70 -345
rect 3 -349 19 -345
rect 6 -353 10 -349
rect 6 -357 40 -353
rect -66 -376 -63 -359
rect -28 -361 -12 -360
rect -28 -365 -16 -361
rect -290 -384 -70 -381
rect -290 -394 -88 -390
rect -284 -403 -280 -394
rect -239 -403 -235 -394
rect -176 -400 -171 -394
rect -137 -400 -132 -394
rect -272 -443 -271 -403
rect -263 -443 -262 -403
rect -276 -448 -258 -443
rect -227 -443 -226 -403
rect -218 -443 -217 -403
rect -254 -452 -250 -443
rect -231 -448 -213 -443
rect -172 -420 -171 -400
rect -133 -420 -132 -400
rect -120 -402 -116 -394
rect -104 -402 -100 -394
rect -185 -429 -180 -420
rect -185 -433 -167 -429
rect -146 -430 -141 -420
rect -112 -430 -108 -422
rect -96 -430 -92 -422
rect -146 -433 -119 -430
rect -209 -450 -205 -443
rect -185 -444 -180 -433
rect -146 -444 -141 -433
rect -112 -433 -103 -430
rect -112 -443 -108 -433
rect -96 -434 -87 -430
rect -96 -443 -92 -434
rect -290 -456 -283 -452
rect -254 -456 -238 -452
rect -284 -473 -280 -469
rect -254 -467 -250 -456
rect -271 -469 -250 -467
rect -276 -470 -250 -469
rect -239 -473 -235 -469
rect -209 -467 -205 -455
rect -226 -469 -205 -467
rect -231 -470 -205 -469
rect -193 -467 -189 -464
rect -176 -467 -172 -464
rect -193 -470 -172 -467
rect -168 -473 -163 -464
rect -154 -467 -150 -464
rect -137 -467 -133 -464
rect -154 -470 -133 -467
rect -129 -473 -124 -464
rect -120 -473 -116 -447
rect -104 -473 -100 -447
rect -74 -473 -70 -384
rect -67 -379 -63 -376
rect -67 -390 -64 -379
rect -56 -387 -46 -382
rect 0 -370 4 -365
rect 27 -373 35 -369
rect -67 -393 -63 -390
rect -66 -396 -63 -393
rect -66 -400 -50 -396
rect -58 -468 -55 -400
rect -38 -404 -34 -388
rect -8 -389 -4 -381
rect 0 -381 7 -377
rect 0 -389 3 -381
rect -19 -393 -15 -389
rect -8 -393 3 -389
rect -8 -396 -4 -393
rect 0 -395 3 -393
rect 31 -389 35 -373
rect 0 -399 17 -395
rect -16 -410 -12 -406
rect -34 -414 -13 -410
rect -52 -418 -42 -414
rect 0 -415 4 -399
rect 31 -403 35 -394
rect 10 -410 14 -406
rect 27 -407 35 -403
rect 1 -418 4 -415
rect -52 -453 -47 -418
rect 1 -421 32 -418
rect -28 -424 -2 -421
rect -5 -427 29 -424
rect -16 -432 -8 -429
rect -39 -441 -35 -437
rect -12 -438 -8 -432
rect 25 -437 29 -427
rect 21 -441 29 -437
rect -15 -449 1 -445
rect -12 -452 -8 -449
rect -52 -457 -35 -453
rect -7 -457 1 -453
rect -290 -477 -70 -473
rect -52 -477 -47 -457
rect -39 -465 -35 -461
rect 25 -461 29 -441
rect -12 -468 -8 -464
rect 21 -465 29 -461
rect 33 -462 36 -422
rect -21 -471 -8 -468
rect -290 -478 -47 -477
rect -74 -482 -25 -478
rect 25 -478 29 -465
rect 21 -482 29 -478
rect -15 -490 1 -486
rect -12 -494 -8 -490
rect -12 -498 27 -494
rect 23 -501 27 -498
rect 33 -506 36 -467
rect 41 -471 45 -358
rect 51 -379 54 -289
rect 58 -367 62 -225
rect 68 -259 71 -139
rect 77 -164 81 -76
rect 87 -81 90 -12
rect 101 -35 105 -27
rect 109 -28 113 -27
rect 129 -10 150 -7
rect 129 -11 146 -10
rect 138 -21 142 -11
rect 158 -17 161 -7
rect 220 -5 224 0
rect 290 3 294 19
rect 322 23 325 25
rect 329 23 333 26
rect 322 19 333 23
rect 340 19 344 23
rect 322 11 325 19
rect 318 7 325 11
rect 329 11 333 19
rect 359 18 363 34
rect 290 -1 298 3
rect 240 -9 252 -5
rect 236 -10 252 -9
rect 266 -10 270 -2
rect 321 -5 325 0
rect 341 -9 353 -5
rect 337 -10 353 -9
rect 271 -13 274 -12
rect 367 -13 371 -2
rect 271 -14 276 -13
rect 354 -14 371 -13
rect 271 -17 371 -14
rect 379 -16 383 49
rect 404 59 408 68
rect 449 59 453 68
rect 512 62 517 68
rect 551 62 556 68
rect 416 19 417 59
rect 425 19 426 59
rect 400 10 401 15
rect 412 14 430 19
rect 461 19 462 59
rect 470 19 471 59
rect 434 10 438 19
rect 457 14 475 19
rect 516 42 517 62
rect 555 42 556 62
rect 568 60 572 68
rect 584 60 588 68
rect 503 33 508 42
rect 503 29 521 33
rect 542 32 547 42
rect 576 32 580 40
rect 592 32 596 40
rect 542 29 569 32
rect 479 12 483 19
rect 503 18 508 29
rect 542 18 547 29
rect 576 29 585 32
rect 576 19 580 29
rect 592 28 602 32
rect 592 19 596 28
rect 400 9 405 10
rect 394 6 405 9
rect 434 6 450 10
rect 404 -11 408 -7
rect 434 -5 438 6
rect 417 -7 438 -5
rect 412 -8 438 -7
rect 449 -11 453 -7
rect 479 -5 483 7
rect 462 -7 483 -5
rect 457 -8 483 -7
rect 495 -5 499 -2
rect 512 -5 516 -2
rect 495 -8 516 -5
rect 520 -11 525 -2
rect 534 -5 538 -2
rect 551 -5 555 -2
rect 534 -8 555 -5
rect 559 -11 564 -2
rect 568 -11 572 15
rect 584 -11 588 15
rect 388 -16 602 -11
rect 158 -21 160 -17
rect 117 -28 121 -27
rect 109 -31 121 -28
rect 153 -23 160 -21
rect 433 -22 655 -19
rect 171 -23 655 -22
rect 153 -24 161 -23
rect 153 -31 156 -24
rect 171 -25 454 -23
rect 171 -26 437 -25
rect 171 -27 174 -26
rect 146 -35 156 -31
rect 161 -30 174 -27
rect 185 -30 189 -26
rect 209 -30 213 -26
rect 95 -40 150 -35
rect 93 -48 99 -44
rect 161 -44 165 -30
rect 105 -48 165 -44
rect 99 -52 103 -48
rect 123 -52 127 -48
rect 107 -81 111 -72
rect 143 -52 147 -48
rect 115 -80 119 -72
rect 87 -85 100 -81
rect 107 -85 114 -81
rect 126 -85 133 -81
rect 151 -81 155 -72
rect 193 -79 197 -70
rect 201 -78 205 -70
rect 178 -80 186 -79
rect 175 -81 186 -80
rect 151 -83 186 -81
rect 193 -83 200 -79
rect 222 -78 226 -70
rect 212 -83 214 -79
rect 245 -50 249 -26
rect 279 -30 283 -26
rect 303 -30 307 -26
rect 230 -79 234 -70
rect 253 -75 257 -70
rect 261 -75 264 -47
rect 253 -78 264 -75
rect 230 -83 246 -79
rect 151 -84 178 -83
rect 151 -85 161 -84
rect 87 -169 90 -85
rect 107 -88 111 -85
rect 130 -86 133 -85
rect 99 -112 103 -108
rect 115 -120 119 -108
rect 151 -88 155 -85
rect 230 -86 234 -83
rect 253 -86 257 -78
rect 287 -79 291 -70
rect 295 -78 299 -70
rect 287 -83 294 -79
rect 316 -78 320 -70
rect 306 -83 308 -79
rect 339 -50 343 -26
rect 373 -30 377 -26
rect 397 -30 401 -26
rect 324 -79 328 -70
rect 324 -83 340 -79
rect 324 -86 328 -83
rect 347 -86 351 -70
rect 381 -79 385 -70
rect 389 -78 393 -70
rect 367 -83 374 -79
rect 381 -83 388 -79
rect 410 -78 414 -70
rect 400 -83 402 -79
rect 433 -50 437 -26
rect 457 -32 461 -23
rect 502 -32 506 -23
rect 565 -29 570 -23
rect 604 -29 609 -23
rect 418 -79 422 -70
rect 441 -79 445 -70
rect 469 -72 470 -32
rect 478 -72 479 -32
rect 465 -77 483 -72
rect 514 -72 515 -32
rect 523 -72 524 -32
rect 418 -83 434 -79
rect 441 -81 454 -79
rect 487 -81 491 -72
rect 510 -77 528 -72
rect 569 -49 570 -29
rect 608 -49 609 -29
rect 621 -31 625 -23
rect 637 -31 641 -23
rect 556 -58 561 -49
rect 556 -62 574 -58
rect 595 -59 600 -49
rect 629 -59 633 -51
rect 645 -59 649 -51
rect 595 -62 622 -59
rect 532 -79 536 -72
rect 556 -73 561 -62
rect 595 -73 600 -62
rect 629 -62 638 -59
rect 629 -72 633 -62
rect 645 -63 655 -59
rect 645 -72 649 -63
rect 441 -83 458 -81
rect 418 -86 422 -83
rect 441 -86 445 -83
rect 451 -85 458 -83
rect 487 -85 503 -81
rect 123 -112 127 -108
rect 143 -114 147 -98
rect 143 -118 160 -114
rect 185 -114 189 -106
rect 193 -107 197 -106
rect 213 -89 234 -86
rect 213 -90 229 -89
rect 222 -100 226 -90
rect 201 -107 205 -106
rect 193 -110 205 -107
rect 230 -114 234 -110
rect 245 -114 249 -96
rect 279 -114 283 -106
rect 287 -107 291 -106
rect 307 -89 328 -86
rect 307 -90 323 -89
rect 316 -100 320 -90
rect 295 -107 299 -106
rect 287 -110 299 -107
rect 324 -114 328 -110
rect 339 -114 343 -96
rect 373 -114 377 -106
rect 381 -107 385 -106
rect 401 -89 422 -86
rect 401 -90 417 -89
rect 410 -100 414 -90
rect 389 -107 393 -106
rect 381 -110 393 -107
rect 418 -114 422 -110
rect 433 -102 437 -96
rect 457 -102 461 -98
rect 487 -96 491 -85
rect 470 -98 491 -96
rect 465 -99 491 -98
rect 502 -102 506 -98
rect 532 -96 536 -84
rect 515 -98 536 -96
rect 510 -99 536 -98
rect 548 -96 552 -93
rect 565 -96 569 -93
rect 548 -99 569 -96
rect 573 -102 578 -93
rect 587 -96 591 -93
rect 604 -96 608 -93
rect 587 -99 608 -96
rect 612 -102 617 -93
rect 621 -102 625 -76
rect 637 -102 641 -76
rect 433 -107 655 -102
rect 433 -114 437 -107
rect 165 -118 394 -114
rect 143 -119 394 -118
rect 143 -120 147 -119
rect 400 -119 437 -114
rect 443 -111 447 -107
rect 115 -125 147 -120
rect 451 -111 477 -110
rect 456 -113 477 -111
rect 473 -124 477 -113
rect 488 -111 492 -107
rect 496 -111 522 -110
rect 501 -113 522 -111
rect 93 -136 98 -132
rect 186 -132 326 -128
rect 437 -125 444 -124
rect 437 -128 439 -125
rect 103 -136 190 -132
rect 210 -136 214 -132
rect 234 -136 238 -132
rect 99 -140 103 -136
rect 118 -140 122 -136
rect 137 -140 141 -136
rect 156 -140 160 -136
rect 172 -140 176 -136
rect 107 -163 111 -160
rect 126 -163 130 -160
rect 145 -163 149 -160
rect 164 -163 168 -160
rect 107 -166 168 -163
rect 164 -167 168 -166
rect 180 -167 184 -160
rect 68 -268 71 -264
rect 77 -342 81 -169
rect 87 -173 100 -169
rect 87 -248 90 -173
rect 164 -171 173 -167
rect 180 -171 189 -167
rect 164 -177 168 -171
rect 180 -174 184 -171
rect 218 -165 222 -156
rect 255 -136 259 -132
rect 226 -164 230 -156
rect 218 -169 225 -165
rect 243 -165 247 -147
rect 341 -145 344 -129
rect 473 -128 489 -124
rect 518 -125 522 -113
rect 534 -113 555 -110
rect 534 -116 538 -113
rect 551 -116 555 -113
rect 451 -137 469 -132
rect 237 -169 247 -165
rect 263 -165 267 -156
rect 314 -159 319 -145
rect 341 -151 345 -145
rect 338 -155 354 -151
rect 319 -163 328 -159
rect 398 -159 402 -143
rect 374 -163 402 -159
rect 263 -169 271 -165
rect 218 -172 222 -169
rect 263 -172 267 -169
rect 99 -223 103 -217
rect 107 -220 122 -217
rect 126 -220 141 -217
rect 172 -204 176 -184
rect 210 -196 214 -192
rect 226 -204 230 -192
rect 234 -196 238 -192
rect 314 -181 319 -165
rect 255 -194 259 -182
rect 314 -185 328 -181
rect 314 -194 319 -185
rect 349 -185 354 -181
rect 349 -186 394 -185
rect 349 -192 354 -186
rect 255 -200 319 -194
rect 349 -193 394 -192
rect 349 -197 354 -193
rect 255 -204 259 -200
rect 314 -201 319 -200
rect 172 -209 273 -204
rect 314 -206 328 -201
rect 398 -201 402 -163
rect 455 -177 456 -137
rect 464 -177 465 -137
rect 473 -137 477 -128
rect 496 -137 514 -132
rect 500 -177 501 -137
rect 509 -177 510 -137
rect 518 -137 522 -130
rect 559 -116 564 -107
rect 573 -113 594 -110
rect 573 -116 577 -113
rect 590 -116 594 -113
rect 598 -116 603 -107
rect 607 -133 611 -107
rect 623 -133 627 -107
rect 542 -147 547 -136
rect 581 -147 586 -136
rect 542 -151 560 -147
rect 542 -160 547 -151
rect 581 -150 608 -147
rect 615 -147 619 -137
rect 631 -146 635 -137
rect 615 -150 624 -147
rect 631 -150 641 -146
rect 581 -160 586 -150
rect 615 -158 619 -150
rect 631 -158 635 -150
rect 443 -186 447 -177
rect 488 -186 492 -177
rect 555 -180 556 -160
rect 594 -180 595 -160
rect 551 -186 556 -180
rect 590 -186 595 -180
rect 607 -186 611 -178
rect 623 -186 627 -178
rect 437 -190 641 -186
rect 145 -220 160 -217
rect 172 -223 176 -209
rect 314 -211 319 -206
rect 394 -205 402 -201
rect 99 -227 176 -223
rect 111 -228 176 -227
rect 194 -216 292 -212
rect 101 -235 103 -231
rect 194 -231 198 -216
rect 108 -235 198 -231
rect 210 -220 214 -216
rect 234 -220 238 -216
rect 257 -220 261 -216
rect 107 -239 111 -235
rect 126 -239 130 -235
rect 145 -239 149 -235
rect 164 -239 168 -235
rect 180 -239 184 -235
rect 218 -249 222 -240
rect 274 -220 278 -216
rect 315 -223 319 -211
rect 226 -248 230 -240
rect 249 -248 253 -240
rect 218 -253 225 -249
rect 237 -253 244 -249
rect 260 -253 267 -249
rect 282 -249 286 -240
rect 315 -237 320 -223
rect 341 -229 345 -223
rect 338 -233 354 -229
rect 315 -241 328 -237
rect 398 -237 402 -205
rect 440 -203 444 -190
rect 440 -207 453 -203
rect 505 -204 506 -197
rect 523 -203 528 -197
rect 374 -241 422 -237
rect 282 -253 291 -249
rect 218 -256 222 -253
rect 115 -262 119 -259
rect 134 -262 138 -259
rect 153 -262 157 -259
rect 172 -262 176 -259
rect 115 -265 176 -262
rect 172 -266 176 -265
rect 188 -266 192 -259
rect 172 -270 181 -266
rect 188 -270 195 -266
rect 172 -276 176 -270
rect 188 -273 192 -270
rect 107 -322 111 -316
rect 115 -319 130 -316
rect 134 -319 149 -316
rect 180 -298 184 -283
rect 210 -290 214 -286
rect 226 -290 230 -286
rect 241 -259 244 -253
rect 234 -290 238 -286
rect 249 -298 253 -286
rect 264 -275 267 -253
rect 282 -256 286 -253
rect 315 -258 320 -241
rect 315 -262 328 -258
rect 257 -290 261 -286
rect 274 -298 278 -266
rect 315 -279 320 -262
rect 349 -262 354 -258
rect 349 -263 414 -262
rect 349 -270 354 -263
rect 349 -271 414 -270
rect 349 -275 354 -271
rect 315 -284 328 -279
rect 315 -297 320 -284
rect 349 -283 354 -279
rect 349 -284 414 -283
rect 349 -291 354 -284
rect 349 -292 414 -291
rect 349 -296 354 -292
rect 289 -298 320 -297
rect 180 -300 320 -298
rect 180 -303 328 -300
rect 153 -319 168 -316
rect 180 -322 184 -303
rect 315 -305 328 -303
rect 418 -300 422 -241
rect 107 -327 184 -322
rect 189 -310 297 -306
rect 105 -335 114 -331
rect 189 -331 193 -310
rect 119 -335 193 -331
rect 210 -314 214 -310
rect 234 -314 238 -310
rect 259 -314 263 -310
rect 111 -339 115 -335
rect 135 -339 139 -335
rect 158 -339 162 -335
rect 119 -368 123 -359
rect 175 -339 179 -335
rect 218 -343 222 -334
rect 279 -314 283 -310
rect 321 -328 327 -305
rect 414 -304 422 -300
rect 226 -342 230 -334
rect 251 -342 255 -334
rect 218 -347 225 -343
rect 237 -345 246 -343
rect 237 -347 241 -345
rect 218 -350 222 -347
rect 262 -345 269 -343
rect 262 -347 266 -345
rect 287 -343 291 -334
rect 315 -332 327 -328
rect 287 -347 296 -343
rect 315 -345 320 -332
rect 343 -337 347 -331
rect 340 -341 356 -337
rect 287 -350 291 -347
rect 127 -367 131 -359
rect 150 -367 154 -359
rect 98 -372 112 -368
rect 119 -372 126 -368
rect 138 -372 145 -368
rect 161 -372 168 -368
rect 183 -368 187 -359
rect 183 -372 193 -368
rect 51 -444 54 -384
rect 58 -435 62 -372
rect 119 -375 123 -372
rect 111 -409 115 -405
rect 127 -409 131 -405
rect 142 -378 145 -372
rect 135 -409 139 -405
rect 150 -417 154 -405
rect 165 -394 168 -372
rect 183 -375 187 -372
rect 210 -384 214 -380
rect 226 -384 230 -380
rect 175 -391 179 -385
rect 234 -384 238 -380
rect 175 -392 204 -391
rect 251 -392 255 -380
rect 259 -384 263 -380
rect 315 -349 330 -345
rect 418 -345 422 -304
rect 440 -248 444 -207
rect 519 -207 528 -203
rect 493 -215 498 -211
rect 453 -216 498 -215
rect 519 -216 520 -211
rect 493 -224 498 -216
rect 453 -225 498 -224
rect 493 -229 498 -225
rect 517 -233 520 -216
rect 493 -237 520 -233
rect 440 -252 453 -248
rect 502 -249 506 -237
rect 523 -248 528 -207
rect 440 -311 444 -252
rect 519 -252 528 -248
rect 493 -260 498 -256
rect 453 -261 498 -260
rect 519 -261 520 -256
rect 493 -269 498 -261
rect 453 -270 498 -269
rect 493 -274 498 -270
rect 517 -278 520 -261
rect 493 -282 500 -278
rect 505 -282 520 -278
rect 514 -298 520 -294
rect 470 -307 494 -302
rect 440 -315 450 -311
rect 440 -316 470 -315
rect 440 -345 444 -316
rect 479 -320 483 -307
rect 517 -311 520 -298
rect 514 -315 520 -311
rect 523 -319 528 -252
rect 514 -324 528 -319
rect 514 -337 520 -333
rect 376 -349 444 -345
rect 470 -346 494 -341
rect 279 -363 283 -360
rect 315 -363 320 -349
rect 440 -350 444 -349
rect 440 -354 450 -350
rect 440 -355 470 -354
rect 279 -367 320 -363
rect 279 -368 330 -367
rect 279 -392 283 -368
rect 175 -397 283 -392
rect 315 -371 330 -368
rect 440 -367 444 -355
rect 315 -389 320 -371
rect 351 -371 356 -367
rect 351 -372 436 -371
rect 440 -371 452 -367
rect 480 -368 483 -346
rect 517 -350 520 -337
rect 514 -354 520 -350
rect 523 -358 528 -324
rect 514 -363 528 -358
rect 523 -367 528 -363
rect 351 -380 356 -372
rect 351 -381 436 -380
rect 351 -385 356 -381
rect 440 -383 444 -371
rect 497 -371 528 -367
rect 472 -379 493 -375
rect 440 -387 452 -383
rect 480 -384 483 -379
rect 523 -383 528 -371
rect 315 -394 330 -389
rect 158 -409 162 -405
rect 175 -417 179 -397
rect 105 -421 179 -417
rect 200 -404 269 -400
rect 110 -422 178 -421
rect 200 -425 203 -404
rect 107 -429 203 -425
rect 210 -408 214 -404
rect 234 -408 238 -404
rect 104 -433 108 -429
rect 128 -433 132 -429
rect 112 -462 116 -453
rect 145 -433 149 -429
rect 218 -437 222 -428
rect 251 -408 255 -404
rect 226 -436 230 -428
rect 218 -441 225 -437
rect 237 -441 244 -437
rect 259 -437 263 -428
rect 315 -411 320 -394
rect 351 -393 356 -389
rect 351 -394 436 -393
rect 351 -402 356 -394
rect 351 -403 436 -402
rect 351 -407 356 -403
rect 315 -416 330 -411
rect 315 -432 320 -416
rect 351 -415 356 -411
rect 351 -416 436 -415
rect 351 -423 356 -416
rect 351 -424 436 -423
rect 351 -428 356 -424
rect 259 -441 266 -437
rect 315 -437 330 -432
rect 440 -432 444 -387
rect 497 -387 528 -383
rect 472 -395 493 -391
rect 480 -401 484 -395
rect 218 -444 222 -441
rect 120 -461 124 -453
rect 98 -466 105 -462
rect 112 -466 119 -462
rect 131 -466 138 -462
rect 153 -462 157 -453
rect 153 -466 163 -462
rect 112 -469 116 -466
rect 104 -493 108 -489
rect 120 -501 124 -489
rect 135 -470 138 -466
rect 153 -469 157 -466
rect 210 -468 214 -464
rect 128 -493 132 -489
rect 226 -476 230 -464
rect 241 -445 244 -441
rect 259 -444 263 -441
rect 234 -468 238 -464
rect 315 -443 320 -437
rect 436 -436 444 -432
rect 524 -443 528 -387
rect 315 -446 528 -443
rect 251 -476 255 -454
rect 315 -476 320 -446
rect 145 -482 149 -479
rect 204 -481 320 -476
rect 190 -482 209 -481
rect 145 -488 209 -482
rect 145 -501 149 -488
rect 120 -506 149 -501
<< m2contact >>
rect 457 94 462 99
<< metal2 >>
rect 219 158 223 159
rect 219 154 388 158
rect -25 140 140 143
rect -162 131 -132 134
rect -137 127 -132 131
rect -83 128 -77 132
rect -176 113 -171 122
rect -204 108 -171 113
rect -82 65 -77 128
rect -25 84 -21 140
rect 61 131 91 134
rect 137 133 140 140
rect 86 127 91 131
rect 168 139 201 143
rect 47 113 52 122
rect 19 108 52 113
rect 168 111 171 139
rect 151 107 171 111
rect 219 106 223 154
rect 321 138 359 141
rect 254 121 255 128
rect 321 106 325 138
rect -25 81 -18 84
rect -21 75 -18 81
rect -25 71 -18 75
rect -82 59 -44 65
rect -162 37 -132 40
rect -137 33 -132 37
rect -82 35 -59 40
rect -176 19 -171 28
rect -204 14 -171 19
rect -162 -57 -132 -54
rect -137 -61 -132 -57
rect -176 -75 -171 -66
rect -204 -80 -171 -75
rect -87 -93 -83 -60
rect -63 -64 -59 35
rect -49 -5 -44 59
rect -25 27 -21 71
rect 184 67 187 96
rect 192 91 242 96
rect 294 91 344 96
rect 355 81 359 138
rect 383 109 387 154
rect 516 126 546 129
rect 541 122 546 126
rect 383 104 388 109
rect 502 108 507 117
rect 393 104 395 106
rect 383 102 395 104
rect 474 103 507 108
rect 355 77 399 81
rect 97 64 187 67
rect 35 29 85 34
rect -25 23 -18 27
rect -12 23 -9 27
rect 33 -4 37 29
rect 46 8 63 13
rect 97 4 100 64
rect 351 62 353 67
rect 351 53 354 62
rect 351 49 366 53
rect 220 34 224 44
rect 321 34 325 47
rect 129 26 182 29
rect 129 5 132 26
rect 179 24 182 26
rect 179 19 188 24
rect 193 19 243 24
rect 294 19 344 24
rect 68 1 100 4
rect -49 -9 33 -5
rect -49 -10 6 -9
rect 10 -38 15 -18
rect 47 -34 52 -29
rect -1 -50 28 -47
rect 48 -51 52 -34
rect 47 -56 52 -51
rect -63 -68 -34 -64
rect -87 -97 -44 -93
rect -47 -146 -44 -97
rect -37 -112 -34 -68
rect 68 -80 71 1
rect 120 0 121 4
rect 130 0 132 5
rect 116 -4 120 -1
rect 137 -4 142 0
rect 116 -7 142 -4
rect 150 -68 153 -18
rect 179 -19 182 19
rect 363 -18 366 49
rect 394 15 399 77
rect 526 30 556 33
rect 551 26 556 30
rect 512 12 517 21
rect 394 6 399 9
rect 484 7 517 12
rect 179 -22 345 -19
rect 78 -71 153 -68
rect 213 -74 216 -22
rect 269 -31 273 -26
rect 269 -51 272 -31
rect 114 -79 144 -75
rect 114 -80 119 -79
rect 68 -83 78 -80
rect 16 -112 66 -107
rect 14 -145 18 -112
rect 75 -121 78 -83
rect 139 -80 144 -79
rect 214 -79 216 -74
rect 268 -54 272 -51
rect 200 -86 226 -83
rect 103 -117 123 -112
rect 132 -121 135 -91
rect 268 -121 271 -54
rect 307 -74 310 -22
rect 342 -41 345 -22
rect 354 -21 367 -18
rect 354 -32 357 -21
rect 342 -44 404 -41
rect 401 -74 404 -44
rect 579 -61 609 -58
rect 604 -65 609 -61
rect 308 -79 310 -74
rect 275 -114 278 -83
rect 294 -86 320 -83
rect 402 -79 404 -74
rect 565 -79 570 -70
rect 388 -86 414 -83
rect 537 -84 570 -79
rect 275 -117 295 -114
rect 66 -122 156 -121
rect 171 -122 246 -121
rect 66 -125 246 -122
rect 268 -124 276 -121
rect 27 -133 44 -128
rect 66 -134 71 -125
rect 132 -126 135 -125
rect 243 -142 246 -125
rect 273 -136 276 -124
rect -162 -150 -132 -147
rect -137 -154 -132 -150
rect -86 -153 -57 -149
rect -47 -150 14 -146
rect 291 -149 294 -117
rect 328 -119 331 -97
rect -176 -168 -171 -159
rect -204 -173 -171 -168
rect -61 -236 -57 -153
rect 275 -152 294 -149
rect 307 -122 331 -119
rect 275 -158 278 -152
rect -9 -179 -4 -159
rect 90 -163 210 -160
rect 90 -164 93 -163
rect 82 -169 93 -164
rect 225 -163 256 -159
rect 275 -161 283 -158
rect 225 -164 230 -163
rect 28 -175 33 -170
rect 251 -164 256 -163
rect -20 -191 9 -188
rect 29 -192 33 -175
rect 28 -197 33 -192
rect 214 -201 234 -196
rect 280 -204 283 -161
rect 307 -212 310 -122
rect 523 -130 556 -125
rect 326 -138 397 -135
rect 551 -139 556 -130
rect 590 -148 595 -144
rect 565 -151 595 -148
rect 325 -172 346 -168
rect 325 -173 328 -172
rect 341 -177 349 -172
rect 323 -192 328 -178
rect 498 -197 506 -192
rect 505 -204 506 -197
rect 307 -213 337 -212
rect 307 -215 344 -213
rect 334 -216 344 -215
rect 340 -218 344 -216
rect 63 -224 307 -220
rect 312 -224 314 -220
rect -162 -244 -132 -241
rect -137 -248 -132 -244
rect -86 -248 -62 -245
rect 226 -247 275 -243
rect -176 -262 -171 -253
rect -204 -267 -171 -262
rect -65 -287 -62 -248
rect -1 -253 49 -248
rect 92 -252 206 -248
rect 225 -248 230 -247
rect 248 -248 253 -247
rect 270 -248 275 -247
rect 323 -249 346 -246
rect -3 -286 1 -253
rect 341 -254 349 -249
rect 96 -257 207 -256
rect 68 -259 207 -257
rect 73 -260 101 -259
rect 204 -260 207 -259
rect 73 -264 75 -260
rect 104 -268 107 -265
rect 204 -264 241 -260
rect 10 -274 27 -269
rect 77 -271 108 -268
rect 54 -280 264 -277
rect -65 -291 -3 -287
rect 214 -295 225 -290
rect 239 -295 257 -290
rect -26 -320 -21 -300
rect 11 -316 16 -311
rect -37 -332 -8 -329
rect 12 -333 16 -316
rect 297 -317 301 -267
rect 323 -270 328 -254
rect -162 -338 -132 -335
rect -137 -342 -132 -338
rect 11 -338 16 -333
rect 42 -320 301 -317
rect -176 -356 -171 -347
rect -204 -361 -171 -356
rect -87 -356 -84 -341
rect 42 -353 45 -320
rect 226 -341 280 -337
rect 82 -347 205 -343
rect 225 -342 230 -341
rect 250 -342 255 -341
rect 275 -342 280 -341
rect 305 -344 308 -289
rect 323 -291 328 -275
rect 301 -347 308 -344
rect 500 -311 505 -283
rect -87 -359 -66 -356
rect 127 -366 176 -362
rect 126 -367 131 -366
rect 63 -372 93 -367
rect 149 -367 154 -366
rect 171 -367 176 -366
rect 55 -383 142 -379
rect 214 -389 225 -384
rect 239 -389 259 -384
rect -19 -394 31 -389
rect -21 -427 -17 -394
rect -8 -415 9 -410
rect 91 -419 94 -396
rect 99 -399 165 -396
rect 115 -414 126 -409
rect 140 -414 158 -409
rect 312 -412 315 -315
rect 491 -316 505 -311
rect 37 -422 94 -419
rect 300 -415 315 -412
rect 325 -354 343 -351
rect 325 -358 328 -354
rect 343 -358 348 -354
rect 479 -350 482 -325
rect 479 -355 486 -350
rect 343 -363 351 -358
rect 325 -380 330 -363
rect 325 -402 330 -385
rect -69 -429 -21 -428
rect -162 -432 -132 -429
rect -137 -436 -132 -432
rect -82 -432 -21 -429
rect 225 -435 252 -431
rect 225 -436 230 -435
rect 63 -440 205 -437
rect 247 -436 252 -435
rect 300 -437 303 -415
rect 325 -423 330 -407
rect 271 -441 303 -437
rect -176 -450 -171 -441
rect -204 -455 -171 -450
rect -44 -461 -39 -441
rect 55 -449 241 -447
rect 50 -450 241 -449
rect -7 -457 -2 -452
rect -55 -473 -26 -470
rect -6 -474 -2 -457
rect 119 -460 146 -456
rect 119 -461 124 -460
rect 37 -466 93 -462
rect 141 -461 146 -460
rect -7 -479 -2 -474
rect 45 -475 135 -472
rect 214 -473 234 -468
rect 108 -498 128 -493
<< m123contact >>
rect 135 167 142 173
rect 159 164 165 170
rect -167 130 -162 135
rect -88 128 -83 133
rect -198 122 -193 127
rect -176 122 -171 127
rect -158 122 -153 127
rect -137 122 -132 127
rect -209 108 -204 113
rect -266 99 -261 104
rect -221 99 -216 104
rect -91 74 -86 79
rect -43 99 -38 104
rect 56 130 61 135
rect 25 122 30 127
rect 47 122 52 127
rect 65 122 70 127
rect 86 122 91 127
rect 135 126 140 133
rect 14 108 19 113
rect 146 107 151 113
rect 201 137 208 143
rect 249 121 254 128
rect 2 99 7 104
rect 218 101 223 106
rect 268 98 273 103
rect 320 101 325 106
rect -167 36 -162 41
rect -89 35 -82 40
rect -198 28 -193 33
rect -176 28 -171 33
rect -158 28 -153 33
rect -137 28 -132 33
rect -209 14 -204 19
rect -266 5 -261 10
rect -221 5 -216 10
rect -92 -22 -86 -15
rect -167 -58 -162 -53
rect -88 -60 -83 -55
rect -198 -66 -193 -61
rect -176 -66 -171 -61
rect -158 -66 -153 -61
rect -137 -66 -132 -61
rect -209 -80 -204 -75
rect -266 -89 -261 -84
rect -221 -89 -216 -84
rect 187 91 192 96
rect 242 91 247 96
rect 289 91 294 96
rect 344 91 349 96
rect 511 125 516 130
rect 480 117 485 122
rect 502 117 507 122
rect 520 117 525 122
rect 541 117 546 122
rect 388 104 393 109
rect 370 98 375 103
rect 469 103 474 108
rect 412 94 417 99
rect 20 58 26 63
rect 53 58 58 63
rect -7 36 -2 41
rect 30 29 35 34
rect 85 29 90 34
rect -18 22 -12 27
rect 4 22 9 27
rect 21 -1 26 4
rect 41 8 46 13
rect 63 8 68 13
rect 219 62 224 67
rect 251 62 257 67
rect 261 58 266 63
rect 321 62 326 67
rect 353 62 359 67
rect 112 53 117 58
rect 363 57 369 62
rect 219 29 224 34
rect 269 26 274 31
rect 320 29 325 34
rect 188 19 193 24
rect 243 19 248 24
rect 289 19 294 24
rect 344 19 349 24
rect 33 -9 38 -4
rect 10 -18 15 -13
rect 42 -34 47 -29
rect 10 -43 15 -38
rect -6 -50 -1 -45
rect 28 -50 33 -45
rect 42 -56 47 -51
rect -91 -113 -86 -108
rect 1 -83 7 -78
rect 34 -83 39 -78
rect 115 -1 120 4
rect 125 0 130 5
rect 137 0 142 5
rect 87 -12 92 -7
rect 149 -18 154 -13
rect 99 -48 105 -43
rect 160 -23 166 -17
rect 220 -10 225 -5
rect 252 -10 257 -5
rect 321 -10 326 -5
rect 353 -10 359 -5
rect 266 -15 271 -10
rect 370 26 375 31
rect 521 29 526 34
rect 490 21 495 26
rect 512 21 517 26
rect 530 21 535 26
rect 551 21 556 26
rect 394 9 400 15
rect 479 7 484 12
rect 422 -2 427 3
rect 467 -2 472 3
rect 383 -16 388 -11
rect 76 -76 81 -71
rect 260 -47 265 -42
rect -26 -105 -21 -100
rect 11 -112 16 -107
rect 66 -112 71 -107
rect -37 -118 -31 -112
rect -15 -119 -10 -114
rect 2 -142 7 -137
rect 114 -85 119 -80
rect 139 -85 144 -80
rect 200 -83 205 -78
rect 209 -79 214 -74
rect 221 -83 226 -78
rect 130 -91 135 -86
rect 98 -117 103 -112
rect 123 -117 128 -112
rect 233 -97 238 -92
rect 160 -118 165 -112
rect 354 -37 359 -32
rect 574 -62 579 -57
rect 543 -70 548 -65
rect 565 -70 570 -65
rect 583 -70 588 -65
rect 604 -70 609 -65
rect 275 -83 280 -78
rect 294 -83 299 -78
rect 303 -79 308 -74
rect 315 -83 320 -78
rect 351 -83 357 -78
rect 362 -84 367 -79
rect 388 -83 393 -78
rect 397 -79 402 -74
rect 409 -83 414 -78
rect 532 -84 537 -79
rect 327 -97 332 -92
rect 421 -97 426 -92
rect 475 -93 480 -88
rect 520 -93 525 -88
rect 22 -133 27 -128
rect 44 -133 49 -128
rect 66 -139 71 -134
rect 98 -136 103 -131
rect 273 -141 278 -136
rect -167 -151 -162 -146
rect -92 -153 -86 -148
rect 14 -150 19 -145
rect 243 -147 248 -142
rect -198 -159 -193 -154
rect -176 -159 -171 -154
rect -158 -159 -153 -154
rect -137 -159 -132 -154
rect -209 -173 -204 -168
rect -266 -182 -261 -177
rect -221 -182 -216 -177
rect -91 -207 -86 -202
rect 394 -120 400 -114
rect 461 -121 466 -116
rect 506 -121 511 -116
rect -9 -159 -4 -154
rect 77 -169 82 -164
rect 210 -165 215 -160
rect 23 -175 28 -170
rect 114 -174 119 -169
rect 133 -174 138 -169
rect 152 -174 157 -169
rect 189 -172 195 -167
rect 225 -169 230 -164
rect 251 -169 256 -164
rect 271 -170 276 -165
rect -9 -184 -4 -179
rect -25 -191 -20 -186
rect 9 -191 14 -186
rect 23 -197 28 -192
rect 209 -201 214 -196
rect 234 -201 239 -196
rect 280 -209 285 -204
rect 340 -129 345 -124
rect 439 -130 444 -125
rect 518 -130 523 -125
rect 320 -138 326 -132
rect 397 -143 404 -135
rect 529 -144 534 -139
rect 551 -144 556 -139
rect 569 -144 574 -139
rect 590 -144 595 -139
rect 560 -152 565 -147
rect 314 -165 319 -159
rect 341 -168 346 -163
rect 323 -178 328 -173
rect 349 -177 354 -172
rect 341 -189 346 -184
rect 323 -197 328 -192
rect 498 -204 505 -197
rect 341 -209 346 -204
rect -16 -224 -10 -219
rect 17 -224 22 -219
rect 58 -225 63 -220
rect 307 -224 312 -219
rect 340 -223 345 -218
rect 509 -226 514 -221
rect -57 -236 -49 -228
rect 103 -235 108 -230
rect -167 -245 -162 -240
rect -92 -248 -86 -242
rect -43 -246 -38 -241
rect 341 -246 346 -241
rect -198 -253 -193 -248
rect -176 -253 -171 -248
rect -158 -253 -153 -248
rect -137 -253 -132 -248
rect -209 -267 -204 -262
rect -266 -276 -261 -271
rect -221 -276 -216 -271
rect -6 -253 -1 -248
rect 49 -253 54 -248
rect 87 -253 92 -248
rect 206 -252 211 -247
rect 225 -253 230 -248
rect 248 -253 253 -248
rect 270 -253 275 -248
rect 291 -253 296 -248
rect -32 -260 -27 -255
rect -15 -283 -10 -278
rect 323 -254 328 -249
rect 68 -264 73 -259
rect 107 -268 112 -263
rect 241 -264 246 -259
rect 5 -274 10 -269
rect 27 -274 32 -269
rect 67 -273 72 -268
rect 122 -273 127 -268
rect 141 -273 146 -268
rect 160 -273 165 -268
rect 195 -271 200 -266
rect 297 -267 302 -262
rect 49 -280 54 -275
rect 264 -280 269 -275
rect -3 -291 2 -286
rect 50 -289 55 -284
rect 209 -295 214 -290
rect 225 -295 230 -290
rect 234 -295 239 -290
rect 257 -295 262 -290
rect -88 -300 -83 -295
rect -26 -300 -21 -295
rect 6 -316 11 -311
rect -26 -325 -21 -320
rect -42 -332 -37 -327
rect -8 -332 -3 -327
rect 349 -255 354 -250
rect 341 -266 346 -261
rect 323 -275 328 -270
rect 509 -271 514 -266
rect -167 -339 -162 -334
rect -89 -341 -84 -336
rect 6 -338 11 -333
rect 305 -289 310 -284
rect -198 -347 -193 -342
rect -176 -347 -171 -342
rect -158 -347 -153 -342
rect -137 -347 -132 -342
rect -209 -361 -204 -356
rect 114 -335 119 -330
rect 77 -347 82 -342
rect 205 -347 211 -341
rect 225 -347 230 -342
rect 241 -350 246 -345
rect 250 -347 255 -342
rect 266 -350 271 -345
rect 275 -347 280 -342
rect 296 -347 301 -342
rect 341 -287 346 -282
rect 500 -283 505 -278
rect 323 -296 328 -291
rect 486 -294 491 -289
rect 341 -308 346 -303
rect 312 -315 317 -310
rect -66 -359 -61 -354
rect 40 -358 45 -353
rect -34 -365 -28 -360
rect -1 -365 4 -360
rect -266 -370 -261 -365
rect -221 -370 -216 -365
rect 58 -372 63 -367
rect 93 -372 98 -367
rect 126 -372 131 -367
rect 149 -372 154 -367
rect 171 -372 176 -367
rect 193 -372 198 -367
rect -61 -387 -56 -382
rect 50 -384 55 -379
rect 142 -383 147 -378
rect 209 -389 214 -384
rect 225 -389 230 -384
rect 234 -389 239 -384
rect 259 -389 264 -384
rect -88 -394 -83 -389
rect -24 -394 -19 -389
rect 31 -394 36 -389
rect -50 -401 -45 -396
rect -33 -424 -28 -419
rect -13 -415 -8 -410
rect 9 -415 14 -410
rect 32 -422 37 -417
rect 94 -399 99 -394
rect 165 -399 170 -394
rect 110 -414 115 -409
rect 126 -414 131 -409
rect 135 -414 140 -409
rect 158 -414 163 -409
rect 486 -316 491 -311
rect 478 -325 483 -320
rect 343 -331 348 -326
rect 343 -354 348 -349
rect 486 -334 491 -329
rect 486 -355 491 -350
rect 325 -363 330 -358
rect 351 -363 356 -358
rect 343 -375 348 -370
rect 325 -385 330 -380
rect 343 -397 348 -392
rect 325 -407 330 -402
rect -167 -433 -162 -428
rect -87 -434 -82 -429
rect -21 -432 -16 -427
rect 98 -429 107 -424
rect -198 -441 -193 -436
rect -176 -441 -171 -436
rect -158 -441 -153 -436
rect -137 -441 -132 -436
rect -44 -441 -39 -436
rect 58 -440 63 -435
rect 205 -441 211 -436
rect 225 -441 230 -436
rect 247 -441 252 -436
rect 266 -441 271 -436
rect 343 -419 348 -414
rect 325 -428 330 -423
rect 343 -440 348 -435
rect -209 -455 -204 -450
rect -266 -464 -261 -459
rect -221 -464 -216 -459
rect 50 -449 55 -444
rect 241 -450 246 -445
rect -12 -457 -7 -452
rect -44 -466 -39 -461
rect -60 -473 -55 -468
rect -26 -473 -21 -468
rect 32 -467 37 -462
rect 93 -467 98 -462
rect 119 -466 124 -461
rect 141 -466 146 -461
rect 163 -466 168 -461
rect -12 -479 -7 -474
rect 40 -476 45 -471
rect 135 -475 140 -470
rect 209 -473 214 -468
rect 234 -473 239 -468
rect 103 -498 108 -493
rect 128 -498 133 -493
rect 22 -506 27 -501
<< metal3 >>
rect 142 167 159 170
rect -198 142 -155 146
rect -198 127 -193 142
rect -158 127 -155 142
rect 25 143 151 146
rect 25 142 68 143
rect 25 127 30 142
rect 65 127 68 142
rect -198 104 -194 122
rect 25 104 29 122
rect 146 113 151 143
rect 159 128 162 164
rect 208 137 523 141
rect 159 123 249 128
rect -290 99 -266 104
rect -261 99 -221 104
rect -216 102 -194 104
rect -67 102 -43 104
rect -216 99 -43 102
rect -38 99 2 104
rect 7 99 29 104
rect -290 10 -287 99
rect 159 80 164 123
rect 480 122 485 137
rect 520 122 523 137
rect 251 98 268 103
rect 353 98 370 103
rect 480 99 484 117
rect -60 78 164 80
rect -86 75 164 78
rect -86 74 -71 75
rect -76 59 -71 74
rect -198 48 -155 52
rect -198 33 -193 48
rect -158 33 -155 48
rect -198 10 -194 28
rect -290 5 -266 10
rect -261 5 -221 10
rect -216 5 -194 10
rect -290 -84 -287 5
rect -77 2 -71 59
rect 26 58 53 63
rect 112 58 118 75
rect 251 67 257 98
rect 224 62 251 67
rect -7 2 -4 36
rect 20 27 26 58
rect 117 55 118 58
rect 286 31 289 96
rect 353 67 359 98
rect 388 94 412 99
rect 417 98 484 99
rect 417 94 494 98
rect 326 62 353 67
rect 363 53 366 57
rect 490 45 494 94
rect 490 41 533 45
rect 9 22 26 27
rect 252 26 269 31
rect 278 28 289 31
rect -77 -1 21 2
rect -77 -2 -18 -1
rect -77 -17 -71 -2
rect 252 -5 258 26
rect 137 -7 161 -6
rect 92 -9 220 -7
rect 92 -10 145 -9
rect 158 -10 220 -9
rect 225 -10 252 -5
rect -86 -22 -71 -17
rect 266 -16 271 -15
rect -198 -46 -155 -42
rect -198 -61 -193 -46
rect -158 -61 -155 -46
rect -198 -84 -194 -66
rect -290 -89 -266 -84
rect -261 -89 -221 -84
rect -216 -89 -194 -84
rect -290 -177 -287 -89
rect -77 -110 -71 -22
rect 278 -23 281 28
rect 353 26 370 31
rect 490 26 495 41
rect 530 26 533 41
rect 7 -83 34 -78
rect -86 -113 -71 -110
rect -198 -139 -155 -135
rect -198 -154 -193 -139
rect -158 -154 -155 -139
rect -77 -139 -71 -113
rect -26 -139 -23 -105
rect 1 -114 7 -83
rect 161 -112 165 -23
rect 273 -26 281 -23
rect -10 -119 7 -114
rect 160 -119 165 -118
rect 172 -35 245 -33
rect 286 -35 289 24
rect 353 -5 359 26
rect 490 3 494 21
rect 398 -2 422 3
rect 427 -2 467 3
rect 472 -2 494 3
rect 172 -36 289 -35
rect 172 -129 176 -36
rect 230 -38 289 -36
rect 326 -10 353 -5
rect 321 -41 324 -10
rect 303 -42 324 -41
rect 265 -44 324 -42
rect 265 -45 316 -44
rect 354 -78 357 -37
rect 234 -125 237 -97
rect 234 -128 340 -125
rect -77 -142 2 -139
rect 133 -132 176 -129
rect -198 -177 -194 -159
rect -290 -182 -266 -177
rect -261 -182 -221 -177
rect -216 -182 -194 -177
rect -290 -271 -287 -182
rect -77 -202 -71 -142
rect 133 -169 136 -132
rect 234 -136 259 -135
rect 152 -138 273 -136
rect 152 -139 239 -138
rect 252 -139 273 -138
rect 152 -169 155 -139
rect 362 -152 366 -84
rect 451 -88 457 -2
rect 543 -50 586 -46
rect 543 -65 548 -50
rect 583 -65 586 -50
rect 543 -88 547 -70
rect 451 -93 475 -88
rect 480 -93 520 -88
rect 525 -93 547 -88
rect 388 -115 394 -114
rect 192 -155 366 -152
rect 192 -167 195 -155
rect -86 -207 -71 -202
rect -198 -233 -155 -229
rect -198 -248 -193 -233
rect -158 -248 -155 -233
rect -198 -271 -194 -253
rect -290 -276 -266 -271
rect -261 -276 -221 -271
rect -216 -276 -194 -271
rect -290 -365 -287 -276
rect -77 -280 -71 -207
rect -10 -224 17 -219
rect -43 -280 -40 -246
rect -16 -255 -10 -224
rect 114 -228 117 -174
rect 133 -228 136 -174
rect 152 -228 155 -174
rect 271 -185 276 -170
rect 314 -166 319 -165
rect 271 -188 341 -185
rect 311 -209 341 -206
rect 280 -216 283 -209
rect 280 -219 294 -216
rect 311 -219 314 -209
rect 422 -215 425 -97
rect 451 -116 457 -93
rect 437 -121 461 -116
rect 466 -121 506 -116
rect 511 -121 533 -116
rect 435 -130 439 -125
rect 529 -139 533 -121
rect 529 -159 534 -144
rect 569 -159 572 -144
rect 529 -163 572 -159
rect 529 -197 536 -163
rect 509 -200 536 -197
rect 367 -218 425 -215
rect 114 -231 125 -228
rect 133 -231 144 -228
rect 152 -231 163 -228
rect -27 -260 -10 -255
rect 122 -268 125 -231
rect 141 -268 144 -231
rect 160 -268 163 -231
rect 291 -248 294 -219
rect 312 -224 314 -219
rect 72 -272 96 -270
rect 72 -273 122 -272
rect 93 -275 127 -273
rect -77 -283 -15 -280
rect 141 -279 144 -273
rect 93 -282 144 -279
rect -77 -297 -71 -283
rect 93 -284 96 -282
rect 55 -287 96 -284
rect 160 -286 163 -273
rect 100 -289 163 -286
rect -83 -300 -71 -297
rect -198 -327 -155 -323
rect -198 -342 -193 -327
rect -158 -342 -155 -327
rect -198 -365 -194 -347
rect -290 -370 -266 -365
rect -261 -370 -221 -365
rect -216 -370 -194 -365
rect -290 -459 -287 -370
rect -77 -391 -71 -300
rect 100 -331 103 -289
rect 100 -334 105 -331
rect -28 -365 -1 -360
rect -83 -394 -71 -391
rect -198 -421 -155 -417
rect -198 -436 -193 -421
rect -158 -436 -155 -421
rect -77 -421 -71 -394
rect -61 -421 -58 -387
rect -34 -396 -28 -365
rect 102 -385 105 -334
rect 195 -354 198 -271
rect 243 -345 246 -264
rect 302 -265 341 -262
rect 266 -345 269 -280
rect 310 -287 341 -284
rect 312 -308 341 -305
rect 312 -310 317 -308
rect 367 -312 370 -218
rect 509 -221 514 -200
rect 509 -266 514 -226
rect 509 -289 514 -271
rect 345 -315 370 -312
rect 467 -294 486 -289
rect 491 -293 514 -289
rect 345 -326 348 -315
rect 467 -329 471 -294
rect 467 -332 486 -329
rect 195 -357 315 -354
rect 312 -370 315 -357
rect 94 -388 105 -385
rect 94 -394 97 -388
rect -45 -401 -28 -396
rect 193 -397 196 -372
rect 312 -373 343 -370
rect 312 -397 343 -394
rect 193 -400 315 -397
rect -77 -424 -33 -421
rect 305 -419 343 -416
rect -198 -459 -194 -441
rect -290 -464 -266 -459
rect -261 -464 -221 -459
rect -216 -464 -194 -459
rect 305 -461 308 -419
rect 168 -464 308 -461
rect 312 -440 343 -437
rect 312 -486 315 -440
rect 39 -489 315 -486
rect 39 -502 43 -489
rect 27 -505 43 -502
<< m234contact >>
rect 220 44 225 49
rect 321 47 326 52
rect 273 -31 278 -26
rect 430 -130 435 -125
rect 498 -192 506 -185
<< metal4 >>
rect 322 52 326 53
rect 220 -124 225 44
rect 322 -111 326 47
rect 380 -106 384 -105
rect 380 -111 407 -106
rect 322 -115 384 -111
rect 404 -115 506 -111
rect 220 -125 437 -124
rect 220 -128 430 -125
rect 435 -130 444 -125
rect 502 -185 506 -115
rect 502 -203 506 -192
rect 98 -429 102 -424
<< m345contact >>
rect 254 121 260 128
rect 107 53 112 58
rect 260 53 265 58
rect 357 53 363 58
rect 93 -48 99 -43
rect 261 -16 266 -11
rect 388 -16 393 -11
rect 388 -120 394 -115
rect 93 -136 98 -131
rect 314 -171 319 -166
rect 95 -235 103 -230
rect 109 -335 114 -330
rect 93 -429 98 -424
<< metal5 >>
rect 107 -30 110 53
rect 257 -11 260 121
rect 265 55 357 58
rect 257 -16 261 -11
rect 266 -16 271 -10
rect 257 -17 260 -16
rect 90 -33 110 -30
rect 90 -48 93 -33
rect 93 -131 96 -48
rect 388 -114 393 -16
rect 388 -115 394 -114
rect 93 -230 96 -136
rect 314 -166 319 -159
rect 388 -166 393 -120
rect 319 -171 393 -166
rect 93 -235 95 -230
rect 93 -331 96 -235
rect 93 -335 109 -331
rect 93 -424 96 -335
rect 98 -429 102 -424
<< labels >>
rlabel metal1 4 -54 5 -53 3 gnd
rlabel metal1 59 -215 59 -215 1 G1
rlabel metal1 69 -215 69 -215 1 P1
rlabel m123contact 43 -355 43 -355 1 G2
rlabel metal1 52 -355 52 -355 1 P2
rlabel metal2 -11 -7 -11 -7 1 b0
rlabel metal1 -10 25 -10 25 1 a0
rlabel metal1 -30 -116 -30 -116 1 a1
rlabel metal2 -32 -148 -32 -148 1 b1
rlabel metal1 -46 -257 -46 -257 1 a2
rlabel metal2 -48 -289 -48 -289 1 b2
rlabel metal2 -64 -431 -64 -431 1 b3
rlabel metal2 323 118 323 118 1 t20
rlabel metal1 449 -81 449 -81 7 t16
rlabel m123contact 353 -81 353 -81 1 t15
rlabel metal1 270 -167 270 -167 1 t2
rlabel metal1 266 -439 266 -439 1 t6
rlabel metal1 343 -226 343 -226 1 t7
rlabel metal1 343 -148 343 -148 1 t3
rlabel metal1 345 -334 345 -334 1 t12
rlabel metal1 294 -345 294 -345 1 t5
rlabel metal1 290 -252 290 -252 7 t4
rlabel metal1 187 -169 187 -169 1 t8
rlabel m123contact 196 -268 196 -268 1 t9
rlabel metal1 190 -370 190 -370 1 t10
rlabel m234contact 222 45 222 45 1 t17
rlabel metal2 221 117 221 117 1 t18
rlabel metal1 160 -465 160 -465 1 t11
rlabel metal1 88 -99 88 -99 8 P0
rlabel metal1 79 -99 79 -99 1 G0
rlabel metal1 159 -83 159 -83 7 t1
rlabel metal1 177 -2 177 -2 1 t13
rlabel metal2 180 20 180 20 1 c0
rlabel metal1 261 -76 261 -76 1 t14
rlabel metal1 -288 -454 -288 -454 3 i13
rlabel metal1 -65 -398 -65 -398 1 a3
rlabel metal1 -288 -360 -288 -360 3 i03
rlabel metal1 -288 -266 -288 -266 3 i12
rlabel metal1 -288 -172 -288 -172 3 i02
rlabel metal1 -286 -79 -286 -79 3 i11
rlabel metal1 -287 15 -287 15 3 i01
rlabel metal1 -65 109 -65 109 1 i00
rlabel metal3 -288 101 -288 101 3 Clk
rlabel metal1 653 -61 653 -61 7 Cout
rlabel metal1 589 126 589 126 1 s1
rlabel metal1 599 30 599 30 1 s3
rlabel metal1 482 -399 482 -399 1 s2
rlabel metal1 637 -148 637 -148 1 s0
rlabel metal3 -24 76 -24 76 1 vdd
rlabel metal1 -287 109 -287 109 3 i10
rlabel m234contact 323 48 323 48 1 t19
rlabel metal1 34 -498 34 -498 1 P3
rlabel metal1 24 -497 24 -497 1 G3
<< end >>
