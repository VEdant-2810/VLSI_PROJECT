* SPICE3 file created from 1bitaddie.ext - technology: scmos

.option scale=0.09u

M1000 nandg_0/m1_30_1# Bi nandg_0/m1_26_n48# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 nandg_0/m1_26_n48# Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=500 ps=450
M1002 nandg_0/m1_30_1# Bi vdd nandg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=1040 ps=676
M1003 nandg_0/m1_30_1# Ai vdd nandg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 inverter_0/out inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 inverter_0/out inverter_0/in vdd inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1006 inverter_1/out Cin gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1007 inverter_1/out Cin vdd inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1008 manch_0/clk inverter_2/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1009 manch_0/clk inverter_2/in vdd inverter_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1010 Con inverter_0/out manch_0/m1_24_n50# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1011 manch_0/m1_24_n50# manch_0/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 Con xorg_1/A Cin Gnd nfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1013 Con manch_0/clk vdd manch_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1014 xorg_0/inverter_0/out Ai gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1015 xorg_0/inverter_0/out Ai vdd xorg_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1016 xorg_0/inverter_1/out Bi gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1017 xorg_0/inverter_1/out Bi vdd xorg_0/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1018 xorg_1/A Bi xorg_0/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1019 xorg_0/m1_26_n95# Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 xorg_1/A xorg_0/inverter_1/out xorg_0/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1021 xorg_0/m1_102_n91# xorg_0/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 xorg_0/m1_25_n11# xorg_0/inverter_0/out vdd xorg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1023 xorg_1/A Bi xorg_0/m1_25_n11# xorg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1024 xorg_0/m1_102_n17# Ai vdd xorg_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1025 xorg_1/A xorg_0/inverter_1/out xorg_0/m1_102_n17# xorg_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 xorg_1/inverter_0/out xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1027 xorg_1/inverter_0/out xorg_1/A vdd xorg_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1028 xorg_1/inverter_1/out inverter_1/out gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1029 xorg_1/inverter_1/out inverter_1/out vdd xorg_1/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1030 sum inverter_1/out xorg_1/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1031 xorg_1/m1_26_n95# xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 sum xorg_1/inverter_1/out xorg_1/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1033 xorg_1/m1_102_n91# xorg_1/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 xorg_1/m1_25_n11# xorg_1/inverter_0/out vdd xorg_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1035 sum inverter_1/out xorg_1/m1_25_n11# xorg_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1036 xorg_1/m1_102_n17# xorg_1/A vdd xorg_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1037 sum xorg_1/inverter_1/out xorg_1/m1_102_n17# xorg_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 Bi ff_0/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1039 Bi ff_0/inverter_0/in vdd ff_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1040 ff_0/m1_25_n37# Bin gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1041 ff_0/m1_63_0# ff_0/m1_25_n37# ff_0/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1042 ff_0/m1_58_n52# inverter_2/in gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 ff_0/inverter_0/in inverter_2/in ff_0/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1044 ff_0/m1_106_n52# ff_0/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 ff_0/m1_19_n10# Bin vdd ff_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1046 ff_0/m1_25_n37# inverter_2/in ff_0/m1_19_n10# ff_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1047 ff_0/m1_63_0# inverter_2/in vdd ff_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1048 ff_0/inverter_0/in ff_0/m1_63_0# vdd ff_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1049 Ai ff_1/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1050 Ai ff_1/inverter_0/in vdd ff_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1051 ff_1/m1_25_n37# Ain gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1052 ff_1/m1_63_0# ff_1/m1_25_n37# ff_1/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1053 ff_1/m1_58_n52# inverter_2/in gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 ff_1/inverter_0/in inverter_2/in ff_1/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1055 ff_1/m1_106_n52# ff_1/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 ff_1/m1_19_n10# Ain vdd ff_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1057 ff_1/m1_25_n37# inverter_2/in ff_1/m1_19_n10# ff_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1058 ff_1/m1_63_0# inverter_2/in vdd ff_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1059 ff_1/inverter_0/in ff_1/m1_63_0# vdd ff_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1060 sumo ff_2/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1061 sumo ff_2/inverter_0/in vdd ff_2/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1062 ff_2/m1_25_n37# sum gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1063 ff_2/m1_63_0# ff_2/m1_25_n37# ff_2/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1064 ff_2/m1_58_n52# inverter_2/in gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 ff_2/inverter_0/in inverter_2/in ff_2/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1066 ff_2/m1_106_n52# ff_2/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 ff_2/m1_19_n10# sum vdd ff_2/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1068 ff_2/m1_25_n37# inverter_2/in ff_2/m1_19_n10# ff_2/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1069 ff_2/m1_63_0# inverter_2/in vdd ff_2/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1070 ff_2/inverter_0/in ff_2/m1_63_0# vdd ff_2/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
C0 inverter_2/in xorg_0/inverter_0/out 1.49fF
C1 Cin Gnd 1.24fF
C2 inverter_2/in Gnd 3.24fF
C4 vdd Gnd 1.70fF
C5 sum Gnd 1.47fF
C6 xorg_1/inverter_0/out Gnd 1.68fF
C7 Bi Gnd 1.53fF
C8 xorg_0/inverter_0/out Gnd 1.68fF
C9 Ai Gnd 2.80fF
C10 Con Gnd 3.03fF
C11 manch_0/clk Gnd 1.66fF
