magic
tech scmos
timestamp 1764760221
<< nwell >>
rect -122 -1 -77 34
rect -19 -1 27 34
rect 87 -1 133 34
rect 191 -1 237 34
rect 298 -1 344 34
rect 402 -1 448 34
rect 503 -18 549 17
<< ntransistor >>
rect -60 -15 -40 -13
rect 44 -15 64 -13
rect 152 -15 172 -13
rect 257 -15 277 -13
rect 365 -15 385 -13
rect 469 -15 489 -13
rect -101 -52 -99 -32
rect 3 -52 5 -32
rect 109 -52 111 -32
rect 213 -52 215 -32
rect 320 -52 322 -32
rect 424 -52 426 -32
rect 525 -42 527 -32
rect -101 -93 -99 -73
rect 3 -93 5 -73
rect 109 -93 111 -73
rect 213 -93 215 -73
rect 320 -93 322 -73
rect 424 -93 426 -73
<< ptransistor >>
rect -101 6 -99 26
rect 3 6 5 26
rect 109 6 111 26
rect 213 6 215 26
rect 320 6 322 26
rect 424 6 426 26
rect 525 -11 527 9
<< ndiffusion >>
rect -60 -13 -40 -10
rect 44 -13 64 -10
rect 152 -13 172 -10
rect 257 -13 277 -10
rect 365 -13 385 -10
rect 469 -13 489 -10
rect -60 -18 -40 -15
rect 44 -18 64 -15
rect 152 -18 172 -15
rect 257 -18 277 -15
rect 365 -18 385 -15
rect 469 -18 489 -15
rect -104 -52 -101 -32
rect -99 -52 -96 -32
rect 0 -52 3 -32
rect 5 -52 8 -32
rect 106 -52 109 -32
rect 111 -52 114 -32
rect 210 -52 213 -32
rect 215 -52 218 -32
rect 317 -52 320 -32
rect 322 -52 325 -32
rect 421 -52 424 -32
rect 426 -52 429 -32
rect 522 -42 525 -32
rect 527 -42 530 -32
rect -104 -93 -101 -73
rect -99 -93 -96 -73
rect 0 -93 3 -73
rect 5 -93 8 -73
rect 106 -93 109 -73
rect 111 -93 114 -73
rect 210 -93 213 -73
rect 215 -93 218 -73
rect 317 -93 320 -73
rect 322 -93 325 -73
rect 421 -93 424 -73
rect 426 -93 429 -73
<< pdiffusion >>
rect -104 6 -101 26
rect -99 6 -96 26
rect 0 6 3 26
rect 5 6 8 26
rect 106 6 109 26
rect 111 6 114 26
rect 210 6 213 26
rect 215 6 218 26
rect 317 6 320 26
rect 322 6 325 26
rect 421 6 424 26
rect 426 6 429 26
rect 522 -11 525 9
rect 527 -11 530 9
<< ndcontact >>
rect -60 -10 -40 1
rect 44 -10 64 1
rect 152 -10 172 1
rect 257 -10 277 1
rect 365 -10 385 1
rect 469 -10 489 1
rect -60 -29 -40 -18
rect 44 -29 64 -18
rect 152 -29 172 -18
rect 257 -29 277 -18
rect 365 -29 385 -18
rect 469 -29 489 -18
rect -115 -52 -104 -32
rect -96 -52 -85 -32
rect -11 -52 0 -32
rect 8 -52 19 -32
rect 95 -52 106 -32
rect 114 -52 125 -32
rect 199 -52 210 -32
rect 218 -52 229 -32
rect 306 -52 317 -32
rect 325 -52 336 -32
rect 410 -52 421 -32
rect 429 -52 440 -32
rect 511 -42 522 -32
rect 530 -42 541 -32
rect -115 -93 -104 -73
rect -96 -93 -85 -73
rect -11 -93 0 -73
rect 8 -93 19 -73
rect 95 -93 106 -73
rect 114 -93 125 -73
rect 199 -93 210 -73
rect 218 -93 229 -73
rect 306 -93 317 -73
rect 325 -93 336 -73
rect 410 -93 421 -73
rect 429 -93 440 -73
<< pdcontact >>
rect -115 6 -104 26
rect -96 6 -85 26
rect -11 6 0 26
rect 8 6 19 26
rect 95 6 106 26
rect 114 6 125 26
rect 199 6 210 26
rect 218 6 229 26
rect 306 6 317 26
rect 325 6 336 26
rect 410 6 421 26
rect 429 6 440 26
rect 511 -11 522 9
rect 530 -11 541 9
<< polysilicon >>
rect -101 26 -99 30
rect 3 26 5 30
rect 109 26 111 30
rect 213 26 215 30
rect 320 26 322 30
rect 424 26 426 30
rect 525 9 527 13
rect -101 -9 -99 6
rect 3 -6 5 6
rect 109 -5 111 6
rect 213 -3 215 6
rect 320 -3 322 6
rect 424 -3 426 6
rect -72 -15 -60 -13
rect -40 -15 -36 -13
rect 31 -15 44 -13
rect 64 -15 68 -13
rect 142 -15 152 -13
rect 172 -15 177 -13
rect 249 -15 257 -13
rect 277 -15 281 -13
rect 355 -15 365 -13
rect 385 -15 389 -13
rect 457 -15 469 -13
rect 489 -15 493 -13
rect -101 -32 -99 -19
rect 3 -32 5 -20
rect 109 -32 111 -21
rect 213 -32 215 -23
rect 320 -32 322 -23
rect 424 -32 426 -23
rect 525 -32 527 -11
rect 525 -46 527 -42
rect -101 -55 -99 -52
rect 3 -55 5 -52
rect 109 -55 111 -52
rect 213 -55 215 -52
rect 320 -55 322 -52
rect 424 -55 426 -52
rect -101 -73 -99 -61
rect 3 -73 5 -61
rect 109 -73 111 -61
rect 213 -73 215 -61
rect 320 -73 322 -61
rect 424 -73 426 -61
rect -101 -97 -99 -93
rect 3 -97 5 -93
rect 109 -97 111 -93
rect 213 -97 215 -93
rect 320 -97 322 -93
rect 424 -97 426 -93
<< polycontact >>
rect 518 -27 525 -20
<< metal1 >>
rect -122 33 497 41
rect -115 26 -104 33
rect -11 26 0 33
rect 95 26 106 33
rect 199 26 210 33
rect 306 26 317 33
rect 410 26 421 33
rect 490 24 497 33
rect 490 16 549 24
rect -96 1 -85 6
rect 8 1 19 6
rect 114 1 125 6
rect 218 1 229 6
rect 325 1 336 6
rect 429 1 440 6
rect 511 9 522 16
rect -96 -10 -60 1
rect 8 -10 44 1
rect 114 -9 152 1
rect 87 -10 152 -9
rect 218 -9 257 1
rect 191 -10 257 -9
rect 325 -9 365 1
rect 298 -10 365 -9
rect 429 -8 469 1
rect 402 -10 469 -8
rect -96 -32 -85 -10
rect -20 -17 19 -10
rect -20 -18 -13 -17
rect -40 -29 -13 -18
rect 8 -32 19 -17
rect 87 -15 125 -10
rect 87 -18 93 -15
rect 64 -29 93 -18
rect 114 -32 125 -15
rect 191 -15 229 -10
rect 191 -18 197 -15
rect 172 -29 197 -18
rect 218 -32 229 -15
rect 298 -15 336 -10
rect 298 -18 305 -15
rect 277 -29 305 -18
rect 325 -32 336 -15
rect 402 -15 440 -10
rect 402 -18 408 -15
rect 385 -29 408 -18
rect 429 -32 440 -15
rect 489 -20 498 -18
rect 530 -20 541 -11
rect 489 -27 518 -20
rect 530 -27 558 -20
rect 489 -29 498 -27
rect 530 -32 541 -27
rect -115 -73 -104 -52
rect -11 -73 0 -52
rect 95 -73 106 -52
rect 199 -73 210 -52
rect 306 -73 317 -52
rect 410 -73 421 -52
rect 530 -59 541 -42
rect 446 -64 541 -59
rect -96 -98 -85 -93
rect 8 -98 19 -93
rect 114 -98 125 -93
rect 218 -98 229 -93
rect 325 -98 336 -93
rect 429 -98 440 -93
rect 446 -98 451 -64
rect 526 -65 541 -64
rect -115 -103 452 -98
<< labels >>
rlabel metal1 556 -23 556 -23 7 Vout
rlabel metal1 160 38 161 39 5 VDD
rlabel metal1 167 -102 167 -102 1 GND
<< end >>
