magic
tech scmos
timestamp 1764782750
<< metal1 >>
rect 27 25 103 29
rect -32 1 0 5
rect -32 -57 -26 1
rect 25 -11 28 1
rect 62 -17 67 25
rect 102 -17 106 1
rect 0 -51 4 -39
rect 27 -41 30 -39
rect 27 -45 50 -41
rect 80 -45 100 -41
rect -62 -62 -24 -57
rect -62 -93 -58 -62
rect 0 -68 4 -56
rect 27 -68 30 -45
rect 100 -60 103 -45
rect 126 -51 130 -45
rect 126 -60 130 -56
rect -62 -97 -52 -93
rect -22 -97 -12 -94
rect -7 -95 3 -94
rect 26 -95 30 -83
rect -7 -97 0 -95
rect -62 -122 -59 -97
rect 65 -108 69 -60
rect 102 -91 106 -79
rect 130 -95 143 -91
rect 100 -108 103 -107
rect 27 -109 103 -108
rect -24 -110 -21 -109
rect 24 -110 103 -109
rect -24 -113 2 -110
rect 27 -112 103 -110
rect 140 -122 143 -95
rect -62 -125 143 -122
<< m2contact >>
rect 130 1 136 6
rect 0 -56 5 -51
rect 126 -56 131 -51
rect -12 -97 -7 -92
<< metal2 >>
rect -12 4 -9 5
rect -12 1 130 4
rect -12 -92 -9 1
rect 5 -56 126 -52
use inverter  inverter_0
timestamp 1764702656
transform -1 0 -32 0 1 -87
box -10 -25 20 18
use nmos  nmos_0
timestamp 1764668464
transform -1 0 20 0 1 -62
box -10 -25 20 -5
use nmos  nmos_1
timestamp 1764668464
transform 1 0 10 0 1 -89
box -10 -25 20 -5
use nmos  nmos_3
timestamp 1764668464
transform -1 0 120 0 1 -85
box -10 -25 20 -5
use nmos  nmos_2
timestamp 1764668464
transform 1 0 110 0 1 -54
box -10 -25 20 -5
use pmos  pmos_1
timestamp 1764668421
transform -1 0 20 0 1 -29
box -10 -11 20 18
use inverter  inverter_1
timestamp 1764702656
transform 1 0 60 0 1 -35
box -10 -25 20 18
use pmos  pmos_3
timestamp 1764668421
transform 1 0 110 0 1 -35
box -10 -11 20 18
use pmos  pmos_0
timestamp 1764668421
transform 1 0 10 0 1 11
box -10 -11 20 18
use pmos  pmos_2
timestamp 1764668421
transform -1 0 120 0 1 11
box -10 -11 20 18
<< labels >>
rlabel metal2 2 3 2 3 3 An
rlabel space 24 -37 24 -37 1 B
rlabel space 4 -97 4 -97 3 A
rlabel metal2 128 3 128 3 7 A
rlabel space 103 -43 103 -43 1 Bn
rlabel space 127 -94 127 -94 7 An
<< end >>
