* SPICE3 file created from mcc_1b.ext - technology: scmos

.option scale=0.09u

.subckt mcc_1b Cc clk P G Coc gnd vdd
M1000 Coc P a_n32_13# Gnd nfet w=6 l=2
+  ad=60 pd=44 as=60 ps=44
M1001 w_n5_n7# G Coc w_n5_n7# nfet w=6 l=2
+  ad=60 pd=44 as=0 ps=0
M1002 w_n5_n7# clk gnd Gnd nfet w=6 l=2
+  ad=0 pd=0 as=30 ps=22
M1003 vdd clk Coc vdd pfet w=6 l=2
+  ad=30 pd=22 as=30 ps=22
M1004 a_n32_13# clk Cc Gnd nfet w=6 l=2
+  ad=0 pd=0 as=30 ps=22
.ends
