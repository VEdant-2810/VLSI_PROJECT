* SPICE3 file created from 1bitaddie.ext - technology: scmos

.include TSMC_180nm.txt
.option scale=0.09u

M1000 nandg_0_m1_30_1 Bi nandg_0_m1_26_n48 Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 nandg_0_m1_26_n48 Ai gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=500 ps=450
M1002 nandg_0_m1_30_1 Bi vdd nandg_0_pmos_0_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=1040 ps=676
M1003 nandg_0_m1_30_1 Ai vdd nandg_0_pmos_1_w_n8_n5 CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 inverter_0_out inverter_0_in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 inverter_0_out inverter_0_in vdd inverter_0_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1006 inverter_1_out Cin gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1007 inverter_1_out Cin vdd inverter_1_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1008 manch_0_clk inverter_2_in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1009 manch_0_clk inverter_2_in vdd inverter_2_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1010 Con inverter_0_out manch_0_m1_24_n50 Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1011 manch_0_m1_24_n50 manch_0_clk gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 Con xorg_1_A Cin Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1013 Con manch_0_clk vdd manch_0_pmos_0_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1014 xorg_0_inverter_0_out Ai gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1015 xorg_0_inverter_0_out Ai vdd xorg_0_inverter_0_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1016 xorg_0_inverter_1_out Bi gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1017 xorg_0_inverter_1_out Bi vdd xorg_0_inverter_1_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1018 xorg_1_A Bi xorg_0_m1_26_n95 Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1019 xorg_0_m1_26_n95 Ai gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 xorg_1_A xorg_0_inverter_1_out xorg_0_m1_102_n91 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1021 xorg_0_m1_102_n91 xorg_0_inverter_0_out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 xorg_0_m1_25_n11 xorg_0_inverter_0_out vdd xorg_0_pmos_0_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1023 xorg_1_A Bi xorg_0_m1_25_n11 xorg_0_pmos_1_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1024 xorg_0_m1_102_n17 Ai vdd xorg_0_pmos_2_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1025 xorg_1_A xorg_0_inverter_1_out xorg_0_m1_102_n17 xorg_0_pmos_3_w_n8_n5 CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 xorg_1_inverter_0_out xorg_1_A gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1027 xorg_1_inverter_0_out xorg_1_A vdd xorg_1_inverter_0_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1028 xorg_1_inverter_1_out inverter_1_out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1029 xorg_1_inverter_1_out inverter_1_out vdd xorg_1_inverter_1_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1030 sum inverter_1_out xorg_1_m1_26_n95 Gnd CMOSN w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1031 xorg_1_m1_26_n95 xorg_1_A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 sum xorg_1_inverter_1_out xorg_1_m1_102_n91 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1033 xorg_1_m1_102_n91 xorg_1_inverter_0_out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 xorg_1_m1_25_n11 xorg_1_inverter_0_out vdd xorg_1_pmos_0_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1035 sum inverter_1_out xorg_1_m1_25_n11 xorg_1_pmos_1_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1036 xorg_1_m1_102_n17 xorg_1_A vdd xorg_1_pmos_2_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1037 sum xorg_1_inverter_1_out xorg_1_m1_102_n17 xorg_1_pmos_3_w_n8_n5 CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 Bi ff_0_inverter_0_in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1039 Bi ff_0_inverter_0_in vdd ff_0_inverter_0_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1040 ff_0_m1_25_n37 Bin gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1041 ff_0_m1_63_0 ff_0_m1_25_n37 ff_0_m1_58_n52 Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1042 ff_0_m1_58_n52 inverter_2_in gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 ff_0_inverter_0_in inverter_2_in ff_0_m1_106_n52 Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1044 ff_0_m1_106_n52 ff_0_m1_63_0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 ff_0_m1_19_n10 Bin vdd ff_0_pmos_0_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1046 ff_0_m1_25_n37 inverter_2_in ff_0_m1_19_n10 ff_0_pmos_1_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1047 ff_0_m1_63_0 inverter_2_in vdd ff_0_pmos_2_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1048 ff_0_inverter_0_in ff_0_m1_63_0 vdd ff_0_pmos_3_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1049 Ai ff_1_inverter_0_in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1050 Ai ff_1_inverter_0_in vdd ff_1_inverter_0_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1051 ff_1_m1_25_n37 Ain gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1052 ff_1_m1_63_0 ff_1_m1_25_n37 ff_1_m1_58_n52 Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1053 ff_1_m1_58_n52 inverter_2_in gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 ff_1_inverter_0_in inverter_2_in ff_1_m1_106_n52 Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1055 ff_1_m1_106_n52 ff_1_m1_63_0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 ff_1_m1_19_n10 Ain vdd ff_1_pmos_0_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1057 ff_1_m1_25_n37 inverter_2_in ff_1_m1_19_n10 ff_1_pmos_1_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1058 ff_1_m1_63_0 inverter_2_in vdd ff_1_pmos_2_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1059 ff_1_inverter_0_in ff_1_m1_63_0 vdd ff_1_pmos_3_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1060 sumo ff_2_inverter_0_in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1061 sumo ff_2_inverter_0_in vdd ff_2_inverter_0_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1062 ff_2_m1_25_n37 sum gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1063 ff_2_m1_63_0 ff_2_m1_25_n37 ff_2_m1_58_n52 Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1064 ff_2_m1_58_n52 inverter_2_in gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 ff_2_inverter_0_in inverter_2_in ff_2_m1_106_n52 Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1066 ff_2_m1_106_n52 ff_2_m1_63_0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 ff_2_m1_19_n10 sum vdd ff_2_pmos_0_w_n8_n5 CMOSP w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1068 ff_2_m1_25_n37 inverter_2_in ff_2_m1_19_n10 ff_2_pmos_1_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1069 ff_2_m1_63_0 inverter_2_in vdd ff_2_pmos_2_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1070 ff_2_inverter_0_in ff_2_m1_63_0 vdd ff_2_pmos_3_w_n8_n5 CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0

Mn1 Coutinv Con gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
Mp1 Coutinv Con vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0

Mn2 Cout Coutinv gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
Mp2 Cout Coutinv vdd vdd CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0



C0 inverter_2_in xorg_0_inverter_0_out 1.49fF
C1 Cin Gnd 1.24fF
C2 inverter_2_in Gnd 3.24fF
C4 vdd Gnd 1.70fF
C5 sum Gnd 1.47fF
C6 xorg_1_inverter_0_out Gnd 1.68fF
C7 Bi Gnd 1.53fF
C8 xorg_0_inverter_0_out Gnd 1.68fF
C9 Ai Gnd 2.80fF
C10 Con Gnd 3.03fF
C11 manch_0_clk Gnd 1.66fF 



*Ai Bi Cin Con Sum Sumo Clk

Vclk clk gnd PULSE(0 1.8 0 100p 100p 25n 50n)
Va Ai 0 PULSE(0 1.8 0 100p 100p 10n 20n)
Vb Bi 0 PULSE(0 1.8 0 100p 100p 20n 40n)
Vc Cin 0 PULSE(0 1.8 0 100p 100p 30n 60n)
Vdd vdd 0 DC 1.8    

.tran 0.1n 200n

.control
run
plot Ai Bi+2 Cin+4 Cout+8 Sum+10 clk+6
.endc   
.end