magic
tech scmos
timestamp 1731358426
<< nwell >>
rect 0 38 65 93
<< ntransistor >>
rect 11 19 13 29
rect 30 19 32 29
rect 52 19 54 29
<< ptransistor >>
rect 11 45 13 85
rect 30 45 32 85
rect 52 45 54 65
<< ndiffusion >>
rect 10 19 11 29
rect 13 19 14 29
rect 29 19 30 29
rect 32 19 33 29
rect 51 19 52 29
rect 54 19 55 29
<< pdiffusion >>
rect 10 45 11 85
rect 13 45 14 85
rect 29 45 30 85
rect 32 45 33 85
rect 51 45 52 65
rect 54 45 55 65
<< ndcontact >>
rect 5 19 10 29
rect 14 19 19 29
rect 25 19 29 29
rect 33 19 38 29
rect 47 19 51 29
rect 55 19 59 29
<< pdcontact >>
rect 6 45 10 85
rect 14 45 18 85
rect 25 45 29 85
rect 33 45 37 85
rect 47 45 51 65
rect 55 45 59 65
<< polysilicon >>
rect 11 85 13 88
rect 30 85 32 88
rect 52 65 54 68
rect 11 29 13 45
rect 30 29 32 45
rect 52 29 54 45
rect 11 16 13 19
rect 30 16 32 19
rect 52 16 54 19
<< polycontact >>
rect 7 32 11 36
rect 26 32 30 36
rect 47 32 52 37
<< metal1 >>
rect 0 89 65 93
rect 6 85 10 89
rect 18 45 19 85
rect 24 45 25 85
rect 14 40 29 45
rect 47 65 51 89
rect 3 32 7 36
rect 22 32 26 36
rect 55 36 59 45
rect 55 32 65 36
rect 55 29 59 32
rect 5 15 10 19
rect 25 15 29 19
rect 47 15 51 19
rect 0 10 65 15
<< metal2 >>
rect 33 37 38 40
rect 33 34 42 37
rect 19 29 33 34
rect 38 32 42 34
<< m123contact >>
rect 33 40 38 45
rect 14 29 19 34
rect 33 29 38 34
rect 42 32 47 37
<< end >>
