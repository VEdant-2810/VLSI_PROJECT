
.include all_subckts.spice

Vdd vdd gnd {SUPPLY}

Vclk clk 0 PULSE(0 {SUPPLY} 2n 100p 100p 30n 60n)
Vd   D   0 PULSE(0 {SUPPLY} 1n 100p 100p 9n 18n)  
*D is delayed by 5ns, for setup time and holdtime violation protection  


Xff1 clk D Q vdd gnd ff_1bit 

Cq Q gnd 10f

.tran 1n 340n 

.control
run

meas tran Q_delay TRIG v(clk) VAL='0.9*V(SUPPLY)' RISE=1 TARG v(Q) VAL='0.9*V(SUPPLY)' RISE=1


plot V(D)+4 V(clk)+2 v(Q)
.endc
.end
