* five bit manchester carry along with flipflop for input and output

.include TSMC_180nm.txt
.param lambda=0.09u
.param SUPPLY=1.8
.param width_N=20*lambda
.global gnd vdd


* -----------------------------------------------------------
* PMOS subcircuit
* Terminals: D G S B
* Parameter: wp (user-specified width)
* -----------------------------------------------------------
.subckt pmos D G S B wp=0

Mp D G S B CMOSP W={wp} L={2*lambda} 
+ AS={5*wp*lambda} PS={10*lambda + 2*wp} 
+ AD={5*wp*lambda} PD={10*lambda + 2*wp}

.ends pmos

* -----------------------------------------------------------
* NMOS subcircuit
* Terminals: D G S B
* Parameter: wn (user-specified width)
* -----------------------------------------------------------
.subckt nmos D G S B wn=0

Mn D G S B CMOSN W={wn} L={2*lambda} 
+ AS={5*wn*lambda} PS={10*lambda + 2*wn} 
+ AD={5*wn*lambda} PD={10*lambda + 2*wn}
.ends nmos

* -----------------------------------------------------------
* 2input XOR subcircuit
* Terminals: A B Y vdd gnd
* -----------------------------------------------------------
.subckt xor2 A B Y vdd gnd

* ===== Inverters to generate A_bar and B_bar =====
* Inverter 1 -> A_bar
C_abar A_BAR gnd 1f
Xpa_invA A_BAR A vdd vdd pmos wp=1.8u
Xna_invA A_BAR A gnd gnd nmos wn=0.9u

* Inverter 2 -> B_bar
C_bbar B_BAR gnd 1f
Xpa_invB B_BAR B vdd vdd pmos wp=1.8u
Xna_invB B_BAR B gnd gnd nmos wn=0.9u

* ===== PTL Pass Network =====
C_yinv Yinv gnd 1f
* Path 1 : Yinv = Abar when B = 0  -> gate = B_BAR, pass A_BAR -> Yinv
Xn1 Yinv B_BAR A_BAR gnd nmos wn=0.9u

* Path 2 : Yinv = A when B = 1 -> gate = B, pass A -> Yinv
Xn2 Yinv B A gnd nmos wn=0.9u

* ===== Output Inverter (restores swing) =====
Xpa_out Y Yinv vdd vdd pmos wp=1.8u
Xna_out Y Yinv gnd gnd nmos wn=0.9u


.ends xor2

* -----------------------------------------------------------
* Flip FLop 
*
* Terminals:
*   clk In Qout vdd gnd
* ----------------------------------------------------------- 
.subckt ff_1bit clk In Qout vdd gnd 

Xm1 W In vdd vdd pmos wp=1.8u
Xm2 A clk W vdd pmos wp=1.8u
Xm3 A In gnd gnd nmos wn=0.9u

Xm4 B clk vdd vdd pmos wp=1.8u
Xm5 Y A B gnd nmos wn=0.9u
Xm6 Y clk gnd gnd nmos wn=0.9u

Xm7 Qinv B vdd vdd pmos wp=1.8u
Xm8 Qinv clk Z gnd nmos wn=0.9u
Xm9 Z B gnd gnd nmos wn=0.9u

Xinvn Qout Qinv gnd gnd nmos wn=0.9u
Xinvp Qout Qinv vdd vdd pmos wp=1.8u

Cqinv Qinv gnd 1f
Ca A gnd 1f
Cb B gnd 1f
Cz Z gnd 1f
Cy Y gnd 1f
Cw W gnd 1f

.ends ff_1bit


* -----------------------------------------------------------
* TRUE Manchester Carry Chain Cell 
*
* Terminals:
*   clk A B Cin Cinbar Cout Coutbar Sum vdd gnd
* ----------------------------------------------------------- 
.subckt mcl clk A B Cin Cinbar Cout Coutbar Sum vdd gnd

* ----- 1. Generate P = A XOR B -----
Cp P gnd 1f
Xxor_AB A B P vdd gnd xor2

*---------Propagate Coutbar = Cinbar when P = 1
* Pass transistor: gate = P, pass Cinbar -> Coutbar
XpassP Coutbar P Cinbar gnd nmos wn=2u


*----------PMOS with clock as input  (precharge style)
XclkPMOS Coutbar clk vdd vdd pmos wp=1.8u


*----------Generate G = AB , putting two nmos in series with gates as A
C_ab AB gnd 1f
XnA Coutbar A AB gnd nmos wn=0.9u
C_bclk Bclk gnd 1f
XnB AB B Bclk gnd nmos wn=0.9u

XclkNMOS Bclk clk gnd gnd nmos wn=0.9u


* ----- 4. Restoring inverter : Coutbar to Cout 
Xcout_p Cout Coutbar vdd vdd pmos wp=1.8u
Xcout_n Cout Coutbar gnd gnd nmos wn=1.8u

*----------Calculate sum = p ^ cin
Xsum P Cin Sum vdd gnd xor2

.ends mcl

* -----------------------------------------------------------
* TRUE Manchester Carry Chain for 5 bit adder 
*
* Terminals:
*   clk A0 B0 A1 B1 A2 B2 A3 B3 A4 B4 Cin Cinbar Cout Coutbar S0 S1 S2 S3 S4 vdd gnd
* ----------------------------------------------------------- 
* for 1bit module  clk A B Cin Cinbar Cout Coutbar Sum vdd gnd mc1

.subckt mca_5bit clk A0 B0 A1 B1 A2 B2 A3 B3 A4 B4 Cin Cinbar Cout Coutbar S0 S1 S2 S3 S4 vdd gnd

*---------bit 0------------
Xbit0 clk A0 B0 Cin Cinbar C0 C0bar S0 vdd gnd mcl
C_c0 C0 gnd 1f
C_c0bar C0bar gnd 1f
C_s0 S0 gnd 1f

*----------bit 1--------------
Xbit1 clk A1 B1 C0 C0bar C1 C1bar S1 vdd gnd mcl
C_c1 C1 gnd 1f
C_c1bar C1bar gnd 1f
C_s1 S1 gnd 1f

*----------bit 2-------------
Xbit2 clk A2 B2 C1 C1bar C2 C2bar S2 vdd gnd mcl
C_c2 C2 gnd 1f
C_c2bar C2bar gnd 1f
C_s2 S2 gnd 1f

*----------bit 3-------------
Xbit3 clk A3 B3 C2 C2bar C3 C3bar S3 vdd gnd mcl
C_c3 C3 gnd 1f
C_c3bar C3bar gnd 1f
C_s3 S3 gnd 1f

*----------bit 4-------------
Xbit4 clk A4 B4 C3 C3bar Cout Coutbar S4 vdd gnd mcl
C_cout Cout gnd 1f
C_coutbar Coutbar gnd 1f
C_s4 S4 gnd 1f

.ends mca_5bit

*---------------------------------------------------------
*                  TESTBENCH
*---------------------------------------------------------