* SPICE3 file created from fulladd.ext - technology: scmos

.option scale=0.09u

M1000 1bitaddie_1/inverter_0/in 1bitaddie_1/Bi 1bitaddie_1/nandg_0/m1_26_n48# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1001 1bitaddie_1/nandg_0/m1_26_n48# 1bitaddie_1/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=2700 ps=2430
M1002 1bitaddie_1/inverter_0/in 1bitaddie_1/Bi vdd 1bitaddie_1/nandg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=5600 ps=3640
M1003 1bitaddie_1/inverter_0/in 1bitaddie_1/Ai vdd 1bitaddie_1/nandg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 1bitaddie_1/inverter_0/out 1bitaddie_1/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 1bitaddie_1/inverter_0/out 1bitaddie_1/inverter_0/in vdd 1bitaddie_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1006 1bitaddie_1/inverter_1/out 1bitaddie_1/Cin gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1007 1bitaddie_1/inverter_1/out 1bitaddie_1/Cin vdd 1bitaddie_1/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1008 1bitaddie_1/manch_0/clk 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1009 1bitaddie_1/manch_0/clk 1bitaddie_4/clk vdd 1bitaddie_1/inverter_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1010 1bitaddie_2/Cin 1bitaddie_1/inverter_0/out 1bitaddie_1/manch_0/m1_24_n50# Gnd nfet w=4 l=2
+  ad=60 pd=54 as=40 ps=36
M1011 1bitaddie_1/manch_0/m1_24_n50# 1bitaddie_1/manch_0/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 1bitaddie_2/Cin 1bitaddie_1/xorg_1/A 1bitaddie_1/Cin Gnd nfet w=4 l=2
+  ad=0 pd=0 as=60 ps=54
M1013 1bitaddie_2/Cin 1bitaddie_1/manch_0/clk vdd 1bitaddie_1/manch_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1014 1bitaddie_1/xorg_0/inverter_0/out 1bitaddie_1/Ai gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1015 1bitaddie_1/xorg_0/inverter_0/out 1bitaddie_1/Ai vdd 1bitaddie_1/xorg_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1016 1bitaddie_1/xorg_0/inverter_1/out 1bitaddie_1/Bi gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1017 1bitaddie_1/xorg_0/inverter_1/out 1bitaddie_1/Bi vdd 1bitaddie_1/xorg_0/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1018 1bitaddie_1/xorg_1/A 1bitaddie_1/Bi 1bitaddie_1/xorg_0/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1019 1bitaddie_1/xorg_0/m1_26_n95# 1bitaddie_1/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 1bitaddie_1/xorg_1/A 1bitaddie_1/xorg_0/inverter_1/out 1bitaddie_1/xorg_0/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1021 1bitaddie_1/xorg_0/m1_102_n91# 1bitaddie_1/xorg_0/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 1bitaddie_1/xorg_0/m1_25_n11# 1bitaddie_1/xorg_0/inverter_0/out vdd 1bitaddie_1/xorg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1023 1bitaddie_1/xorg_1/A 1bitaddie_1/Bi 1bitaddie_1/xorg_0/m1_25_n11# 1bitaddie_1/xorg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1024 1bitaddie_1/xorg_0/m1_102_n17# 1bitaddie_1/Ai vdd 1bitaddie_1/xorg_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1025 1bitaddie_1/xorg_1/A 1bitaddie_1/xorg_0/inverter_1/out 1bitaddie_1/xorg_0/m1_102_n17# 1bitaddie_1/xorg_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 1bitaddie_1/xorg_1/inverter_0/out 1bitaddie_1/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1027 1bitaddie_1/xorg_1/inverter_0/out 1bitaddie_1/xorg_1/A vdd 1bitaddie_1/xorg_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1028 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/inverter_1/out gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1029 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/inverter_1/out vdd 1bitaddie_1/xorg_1/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1030 1bitaddie_1/sum 1bitaddie_1/inverter_1/out 1bitaddie_1/xorg_1/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1031 1bitaddie_1/xorg_1/m1_26_n95# 1bitaddie_1/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 1bitaddie_1/sum 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/xorg_1/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1033 1bitaddie_1/xorg_1/m1_102_n91# 1bitaddie_1/xorg_1/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 1bitaddie_1/xorg_1/m1_25_n11# 1bitaddie_1/xorg_1/inverter_0/out vdd 1bitaddie_1/xorg_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1035 1bitaddie_1/sum 1bitaddie_1/inverter_1/out 1bitaddie_1/xorg_1/m1_25_n11# 1bitaddie_1/xorg_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1036 1bitaddie_1/xorg_1/m1_102_n17# 1bitaddie_1/xorg_1/A vdd 1bitaddie_1/xorg_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1037 1bitaddie_1/sum 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/xorg_1/m1_102_n17# 1bitaddie_1/xorg_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 1bitaddie_1/Bi 1bitaddie_1/ff_0/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1039 1bitaddie_1/Bi 1bitaddie_1/ff_0/inverter_0/in vdd 1bitaddie_1/ff_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1040 1bitaddie_1/ff_0/m1_25_n37# B1 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1041 1bitaddie_1/ff_0/m1_63_0# 1bitaddie_1/ff_0/m1_25_n37# 1bitaddie_1/ff_0/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1042 1bitaddie_1/ff_0/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 1bitaddie_1/ff_0/inverter_0/in 1bitaddie_4/clk 1bitaddie_1/ff_0/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1044 1bitaddie_1/ff_0/m1_106_n52# 1bitaddie_1/ff_0/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 1bitaddie_1/ff_0/m1_19_n10# B1 vdd 1bitaddie_1/ff_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1046 1bitaddie_1/ff_0/m1_25_n37# 1bitaddie_4/clk 1bitaddie_1/ff_0/m1_19_n10# 1bitaddie_1/ff_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1047 1bitaddie_1/ff_0/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_1/ff_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1048 1bitaddie_1/ff_0/inverter_0/in 1bitaddie_1/ff_0/m1_63_0# vdd 1bitaddie_1/ff_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1049 1bitaddie_1/Ai 1bitaddie_1/ff_1/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1050 1bitaddie_1/Ai 1bitaddie_1/ff_1/inverter_0/in vdd 1bitaddie_1/ff_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1051 1bitaddie_1/ff_1/m1_25_n37# A1 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1052 1bitaddie_1/ff_1/m1_63_0# 1bitaddie_1/ff_1/m1_25_n37# 1bitaddie_1/ff_1/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1053 1bitaddie_1/ff_1/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 1bitaddie_1/ff_1/inverter_0/in 1bitaddie_4/clk 1bitaddie_1/ff_1/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1055 1bitaddie_1/ff_1/m1_106_n52# 1bitaddie_1/ff_1/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 1bitaddie_1/ff_1/m1_19_n10# A1 vdd 1bitaddie_1/ff_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1057 1bitaddie_1/ff_1/m1_25_n37# 1bitaddie_4/clk 1bitaddie_1/ff_1/m1_19_n10# 1bitaddie_1/ff_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1058 1bitaddie_1/ff_1/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_1/ff_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1059 1bitaddie_1/ff_1/inverter_0/in 1bitaddie_1/ff_1/m1_63_0# vdd 1bitaddie_1/ff_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1060 s1 1bitaddie_1/ff_2/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1061 s1 1bitaddie_1/ff_2/inverter_0/in vdd 1bitaddie_1/ff_2/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1062 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_1/sum gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1063 1bitaddie_1/ff_2/m1_63_0# 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_1/ff_2/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1064 1bitaddie_1/ff_2/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 1bitaddie_1/ff_2/inverter_0/in 1bitaddie_4/clk 1bitaddie_1/ff_2/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1066 1bitaddie_1/ff_2/m1_106_n52# 1bitaddie_1/ff_2/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 1bitaddie_1/ff_2/m1_19_n10# 1bitaddie_1/sum vdd 1bitaddie_1/ff_2/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1068 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_4/clk 1bitaddie_1/ff_2/m1_19_n10# 1bitaddie_1/ff_2/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1069 1bitaddie_1/ff_2/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_1/ff_2/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1070 1bitaddie_1/ff_2/inverter_0/in 1bitaddie_1/ff_2/m1_63_0# vdd 1bitaddie_1/ff_2/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1071 1bitaddie_2/inverter_0/in 1bitaddie_2/Bi 1bitaddie_2/nandg_0/m1_26_n48# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1072 1bitaddie_2/nandg_0/m1_26_n48# 1bitaddie_2/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 1bitaddie_2/inverter_0/in 1bitaddie_2/Bi vdd 1bitaddie_2/nandg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1074 1bitaddie_2/inverter_0/in 1bitaddie_2/Ai vdd 1bitaddie_2/nandg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 1bitaddie_2/inverter_0/out 1bitaddie_2/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1076 1bitaddie_2/inverter_0/out 1bitaddie_2/inverter_0/in vdd 1bitaddie_2/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1077 1bitaddie_2/inverter_1/out 1bitaddie_2/Cin gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1078 1bitaddie_2/inverter_1/out 1bitaddie_2/Cin vdd 1bitaddie_2/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1079 1bitaddie_2/manch_0/clk 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1080 1bitaddie_2/manch_0/clk 1bitaddie_4/clk vdd 1bitaddie_2/inverter_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1081 1bitaddie_3/Cin 1bitaddie_2/inverter_0/out 1bitaddie_2/manch_0/m1_24_n50# Gnd nfet w=4 l=2
+  ad=60 pd=54 as=40 ps=36
M1082 1bitaddie_2/manch_0/m1_24_n50# 1bitaddie_2/manch_0/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 1bitaddie_3/Cin 1bitaddie_2/xorg_1/A 1bitaddie_2/Cin Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 1bitaddie_3/Cin 1bitaddie_2/manch_0/clk vdd 1bitaddie_2/manch_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1085 1bitaddie_2/xorg_0/inverter_0/out 1bitaddie_2/Ai gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1086 1bitaddie_2/xorg_0/inverter_0/out 1bitaddie_2/Ai vdd 1bitaddie_2/xorg_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1087 1bitaddie_2/xorg_0/inverter_1/out 1bitaddie_2/Bi gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1088 1bitaddie_2/xorg_0/inverter_1/out 1bitaddie_2/Bi vdd 1bitaddie_2/xorg_0/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1089 1bitaddie_2/xorg_1/A 1bitaddie_2/Bi 1bitaddie_2/xorg_0/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1090 1bitaddie_2/xorg_0/m1_26_n95# 1bitaddie_2/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 1bitaddie_2/xorg_1/A 1bitaddie_2/xorg_0/inverter_1/out 1bitaddie_2/xorg_0/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1092 1bitaddie_2/xorg_0/m1_102_n91# 1bitaddie_2/xorg_0/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1093 1bitaddie_2/xorg_0/m1_25_n11# 1bitaddie_2/xorg_0/inverter_0/out vdd 1bitaddie_2/xorg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1094 1bitaddie_2/xorg_1/A 1bitaddie_2/Bi 1bitaddie_2/xorg_0/m1_25_n11# 1bitaddie_2/xorg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1095 1bitaddie_2/xorg_0/m1_102_n17# 1bitaddie_2/Ai vdd 1bitaddie_2/xorg_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1096 1bitaddie_2/xorg_1/A 1bitaddie_2/xorg_0/inverter_1/out 1bitaddie_2/xorg_0/m1_102_n17# 1bitaddie_2/xorg_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1097 1bitaddie_2/xorg_1/inverter_0/out 1bitaddie_2/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1098 1bitaddie_2/xorg_1/inverter_0/out 1bitaddie_2/xorg_1/A vdd 1bitaddie_2/xorg_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1099 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/inverter_1/out gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1100 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/inverter_1/out vdd 1bitaddie_2/xorg_1/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1101 1bitaddie_2/sum 1bitaddie_2/inverter_1/out 1bitaddie_2/xorg_1/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1102 1bitaddie_2/xorg_1/m1_26_n95# 1bitaddie_2/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 1bitaddie_2/sum 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/xorg_1/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1104 1bitaddie_2/xorg_1/m1_102_n91# 1bitaddie_2/xorg_1/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1105 1bitaddie_2/xorg_1/m1_25_n11# 1bitaddie_2/xorg_1/inverter_0/out vdd 1bitaddie_2/xorg_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1106 1bitaddie_2/sum 1bitaddie_2/inverter_1/out 1bitaddie_2/xorg_1/m1_25_n11# 1bitaddie_2/xorg_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1107 1bitaddie_2/xorg_1/m1_102_n17# 1bitaddie_2/xorg_1/A vdd 1bitaddie_2/xorg_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1108 1bitaddie_2/sum 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/xorg_1/m1_102_n17# 1bitaddie_2/xorg_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 1bitaddie_2/Bi 1bitaddie_2/ff_0/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1110 1bitaddie_2/Bi 1bitaddie_2/ff_0/inverter_0/in vdd 1bitaddie_2/ff_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1111 1bitaddie_2/ff_0/m1_25_n37# B2 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1112 1bitaddie_2/ff_0/m1_63_0# 1bitaddie_2/ff_0/m1_25_n37# 1bitaddie_2/ff_0/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1113 1bitaddie_2/ff_0/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1114 1bitaddie_2/ff_0/inverter_0/in 1bitaddie_4/clk 1bitaddie_2/ff_0/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1115 1bitaddie_2/ff_0/m1_106_n52# 1bitaddie_2/ff_0/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 1bitaddie_2/ff_0/m1_19_n10# B2 vdd 1bitaddie_2/ff_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1117 1bitaddie_2/ff_0/m1_25_n37# 1bitaddie_4/clk 1bitaddie_2/ff_0/m1_19_n10# 1bitaddie_2/ff_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1118 1bitaddie_2/ff_0/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_2/ff_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1119 1bitaddie_2/ff_0/inverter_0/in 1bitaddie_2/ff_0/m1_63_0# vdd 1bitaddie_2/ff_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1120 1bitaddie_2/Ai 1bitaddie_2/ff_1/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1121 1bitaddie_2/Ai 1bitaddie_2/ff_1/inverter_0/in vdd 1bitaddie_2/ff_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1122 1bitaddie_2/ff_1/m1_25_n37# A2 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1123 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_2/ff_1/m1_25_n37# 1bitaddie_2/ff_1/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1124 1bitaddie_2/ff_1/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 1bitaddie_2/ff_1/inverter_0/in 1bitaddie_4/clk 1bitaddie_2/ff_1/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1126 1bitaddie_2/ff_1/m1_106_n52# 1bitaddie_2/ff_1/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 1bitaddie_2/ff_1/m1_19_n10# A2 vdd 1bitaddie_2/ff_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1128 1bitaddie_2/ff_1/m1_25_n37# 1bitaddie_4/clk 1bitaddie_2/ff_1/m1_19_n10# 1bitaddie_2/ff_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1129 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_2/ff_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1130 1bitaddie_2/ff_1/inverter_0/in 1bitaddie_2/ff_1/m1_63_0# vdd 1bitaddie_2/ff_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1131 s2 1bitaddie_2/ff_2/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1132 s2 1bitaddie_2/ff_2/inverter_0/in vdd 1bitaddie_2/ff_2/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1133 1bitaddie_2/ff_2/m1_25_n37# 1bitaddie_2/sum gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1134 1bitaddie_2/ff_2/m1_63_0# 1bitaddie_2/ff_2/m1_25_n37# 1bitaddie_2/ff_2/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1135 1bitaddie_2/ff_2/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 1bitaddie_2/ff_2/inverter_0/in 1bitaddie_4/clk 1bitaddie_2/ff_2/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1137 1bitaddie_2/ff_2/m1_106_n52# 1bitaddie_2/ff_2/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 1bitaddie_2/ff_2/m1_19_n10# 1bitaddie_2/sum vdd 1bitaddie_2/ff_2/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1139 1bitaddie_2/ff_2/m1_25_n37# 1bitaddie_4/clk 1bitaddie_2/ff_2/m1_19_n10# 1bitaddie_2/ff_2/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1140 1bitaddie_2/ff_2/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_2/ff_2/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1141 1bitaddie_2/ff_2/inverter_0/in 1bitaddie_2/ff_2/m1_63_0# vdd 1bitaddie_2/ff_2/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1142 1bitaddie_3/inverter_0/in 1bitaddie_3/Bi 1bitaddie_3/nandg_0/m1_26_n48# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1143 1bitaddie_3/nandg_0/m1_26_n48# 1bitaddie_3/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 1bitaddie_3/inverter_0/in 1bitaddie_3/Bi vdd 1bitaddie_3/nandg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1145 1bitaddie_3/inverter_0/in 1bitaddie_3/Ai vdd 1bitaddie_3/nandg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 1bitaddie_3/inverter_0/out 1bitaddie_3/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1147 1bitaddie_3/inverter_0/out 1bitaddie_3/inverter_0/in vdd 1bitaddie_3/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1148 1bitaddie_3/inverter_1/out 1bitaddie_3/Cin gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1149 1bitaddie_3/inverter_1/out 1bitaddie_3/Cin vdd 1bitaddie_3/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1150 1bitaddie_3/manch_0/clk 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1151 1bitaddie_3/manch_0/clk 1bitaddie_4/clk vdd 1bitaddie_3/inverter_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1152 1bitaddie_4/Cin 1bitaddie_3/inverter_0/out 1bitaddie_3/manch_0/m1_24_n50# Gnd nfet w=4 l=2
+  ad=60 pd=54 as=40 ps=36
M1153 1bitaddie_3/manch_0/m1_24_n50# 1bitaddie_3/manch_0/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 1bitaddie_4/Cin 1bitaddie_3/xorg_1/A 1bitaddie_3/Cin Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 1bitaddie_4/Cin 1bitaddie_3/manch_0/clk vdd 1bitaddie_3/manch_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1156 1bitaddie_3/xorg_0/inverter_0/out 1bitaddie_3/Ai gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1157 1bitaddie_3/xorg_0/inverter_0/out 1bitaddie_3/Ai vdd 1bitaddie_3/xorg_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1158 1bitaddie_3/xorg_0/inverter_1/out 1bitaddie_3/Bi gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1159 1bitaddie_3/xorg_0/inverter_1/out 1bitaddie_3/Bi vdd 1bitaddie_3/xorg_0/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1160 1bitaddie_3/xorg_1/A 1bitaddie_3/Bi 1bitaddie_3/xorg_0/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1161 1bitaddie_3/xorg_0/m1_26_n95# 1bitaddie_3/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1162 1bitaddie_3/xorg_1/A 1bitaddie_3/xorg_0/inverter_1/out 1bitaddie_3/xorg_0/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1163 1bitaddie_3/xorg_0/m1_102_n91# 1bitaddie_3/xorg_0/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 1bitaddie_3/xorg_0/m1_25_n11# 1bitaddie_3/xorg_0/inverter_0/out vdd 1bitaddie_3/xorg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1165 1bitaddie_3/xorg_1/A 1bitaddie_3/Bi 1bitaddie_3/xorg_0/m1_25_n11# 1bitaddie_3/xorg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1166 1bitaddie_3/xorg_0/m1_102_n17# 1bitaddie_3/Ai vdd 1bitaddie_3/xorg_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1167 1bitaddie_3/xorg_1/A 1bitaddie_3/xorg_0/inverter_1/out 1bitaddie_3/xorg_0/m1_102_n17# 1bitaddie_3/xorg_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 1bitaddie_3/xorg_1/inverter_0/out 1bitaddie_3/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1169 1bitaddie_3/xorg_1/inverter_0/out 1bitaddie_3/xorg_1/A vdd 1bitaddie_3/xorg_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1170 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/inverter_1/out gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1171 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/inverter_1/out vdd 1bitaddie_3/xorg_1/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1172 1bitaddie_3/sum 1bitaddie_3/inverter_1/out 1bitaddie_3/xorg_1/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1173 1bitaddie_3/xorg_1/m1_26_n95# 1bitaddie_3/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 1bitaddie_3/sum 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/xorg_1/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1175 1bitaddie_3/xorg_1/m1_102_n91# 1bitaddie_3/xorg_1/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 1bitaddie_3/xorg_1/m1_25_n11# 1bitaddie_3/xorg_1/inverter_0/out vdd 1bitaddie_3/xorg_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1177 1bitaddie_3/sum 1bitaddie_3/inverter_1/out 1bitaddie_3/xorg_1/m1_25_n11# 1bitaddie_3/xorg_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1178 1bitaddie_3/xorg_1/m1_102_n17# 1bitaddie_3/xorg_1/A vdd 1bitaddie_3/xorg_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1179 1bitaddie_3/sum 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/xorg_1/m1_102_n17# 1bitaddie_3/xorg_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1180 1bitaddie_3/Bi 1bitaddie_3/ff_0/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1181 1bitaddie_3/Bi 1bitaddie_3/ff_0/inverter_0/in vdd 1bitaddie_3/ff_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1182 1bitaddie_3/ff_0/m1_25_n37# B3 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1183 1bitaddie_3/ff_0/m1_63_0# 1bitaddie_3/ff_0/m1_25_n37# 1bitaddie_3/ff_0/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1184 1bitaddie_3/ff_0/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 1bitaddie_3/ff_0/inverter_0/in 1bitaddie_4/clk 1bitaddie_3/ff_0/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1186 1bitaddie_3/ff_0/m1_106_n52# 1bitaddie_3/ff_0/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 1bitaddie_3/ff_0/m1_19_n10# B3 vdd 1bitaddie_3/ff_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1188 1bitaddie_3/ff_0/m1_25_n37# 1bitaddie_4/clk 1bitaddie_3/ff_0/m1_19_n10# 1bitaddie_3/ff_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1189 1bitaddie_3/ff_0/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_3/ff_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1190 1bitaddie_3/ff_0/inverter_0/in 1bitaddie_3/ff_0/m1_63_0# vdd 1bitaddie_3/ff_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1191 1bitaddie_3/Ai 1bitaddie_3/ff_1/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1192 1bitaddie_3/Ai 1bitaddie_3/ff_1/inverter_0/in vdd 1bitaddie_3/ff_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1193 1bitaddie_3/ff_1/m1_25_n37# A3 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1194 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_3/ff_1/m1_25_n37# 1bitaddie_3/ff_1/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1195 1bitaddie_3/ff_1/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 1bitaddie_3/ff_1/inverter_0/in 1bitaddie_4/clk 1bitaddie_3/ff_1/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1197 1bitaddie_3/ff_1/m1_106_n52# 1bitaddie_3/ff_1/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 1bitaddie_3/ff_1/m1_19_n10# A3 vdd 1bitaddie_3/ff_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1199 1bitaddie_3/ff_1/m1_25_n37# 1bitaddie_4/clk 1bitaddie_3/ff_1/m1_19_n10# 1bitaddie_3/ff_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1200 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_3/ff_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1201 1bitaddie_3/ff_1/inverter_0/in 1bitaddie_3/ff_1/m1_63_0# vdd 1bitaddie_3/ff_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1202 s3 1bitaddie_3/ff_2/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1203 s3 1bitaddie_3/ff_2/inverter_0/in vdd 1bitaddie_3/ff_2/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1204 1bitaddie_3/ff_2/m1_25_n37# 1bitaddie_3/sum gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1205 1bitaddie_3/ff_2/m1_63_0# 1bitaddie_3/ff_2/m1_25_n37# 1bitaddie_3/ff_2/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1206 1bitaddie_3/ff_2/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 1bitaddie_3/ff_2/inverter_0/in 1bitaddie_4/clk 1bitaddie_3/ff_2/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1208 1bitaddie_3/ff_2/m1_106_n52# 1bitaddie_3/ff_2/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 1bitaddie_3/ff_2/m1_19_n10# 1bitaddie_3/sum vdd 1bitaddie_3/ff_2/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1210 1bitaddie_3/ff_2/m1_25_n37# 1bitaddie_4/clk 1bitaddie_3/ff_2/m1_19_n10# 1bitaddie_3/ff_2/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1211 1bitaddie_3/ff_2/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_3/ff_2/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1212 1bitaddie_3/ff_2/inverter_0/in 1bitaddie_3/ff_2/m1_63_0# vdd 1bitaddie_3/ff_2/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1213 inverter_0/out inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=40 pd=36 as=0 ps=0
M1214 inverter_0/out inverter_0/in vdd inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1215 inverter_1/out inverter_1/in gnd Gnd nfet w=4 l=2
+  ad=60 pd=54 as=0 ps=0
M1216 inverter_1/out inverter_1/in vdd inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1217 1bitaddie_4/inverter_0/in 1bitaddie_4/Bi 1bitaddie_4/nandg_0/m1_26_n48# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1218 1bitaddie_4/nandg_0/m1_26_n48# 1bitaddie_4/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 1bitaddie_4/inverter_0/in 1bitaddie_4/Bi vdd 1bitaddie_4/nandg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1220 1bitaddie_4/inverter_0/in 1bitaddie_4/Ai vdd 1bitaddie_4/nandg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 1bitaddie_4/inverter_0/out 1bitaddie_4/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1222 1bitaddie_4/inverter_0/out 1bitaddie_4/inverter_0/in vdd 1bitaddie_4/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1223 1bitaddie_4/inverter_1/out 1bitaddie_4/Cin gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1224 1bitaddie_4/inverter_1/out 1bitaddie_4/Cin vdd 1bitaddie_4/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1225 1bitaddie_4/manch_0/clk 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1226 1bitaddie_4/manch_0/clk 1bitaddie_4/clk vdd 1bitaddie_4/inverter_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1227 inverter_1/out 1bitaddie_4/inverter_0/out 1bitaddie_4/manch_0/m1_24_n50# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1228 1bitaddie_4/manch_0/m1_24_n50# 1bitaddie_4/manch_0/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 inverter_1/out 1bitaddie_4/xorg_1/A 1bitaddie_4/Cin Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 inverter_1/out 1bitaddie_4/manch_0/clk vdd 1bitaddie_4/manch_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 1bitaddie_4/xorg_0/inverter_0/out 1bitaddie_4/Ai gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1232 1bitaddie_4/xorg_0/inverter_0/out 1bitaddie_4/Ai vdd 1bitaddie_4/xorg_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1233 1bitaddie_4/xorg_0/inverter_1/out 1bitaddie_4/Bi gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1234 1bitaddie_4/xorg_0/inverter_1/out 1bitaddie_4/Bi vdd 1bitaddie_4/xorg_0/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1235 1bitaddie_4/xorg_1/A 1bitaddie_4/Bi 1bitaddie_4/xorg_0/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1236 1bitaddie_4/xorg_0/m1_26_n95# 1bitaddie_4/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 1bitaddie_4/xorg_1/A 1bitaddie_4/xorg_0/inverter_1/out 1bitaddie_4/xorg_0/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1238 1bitaddie_4/xorg_0/m1_102_n91# 1bitaddie_4/xorg_0/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 1bitaddie_4/xorg_0/m1_25_n11# 1bitaddie_4/xorg_0/inverter_0/out vdd 1bitaddie_4/xorg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1240 1bitaddie_4/xorg_1/A 1bitaddie_4/Bi 1bitaddie_4/xorg_0/m1_25_n11# 1bitaddie_4/xorg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1241 1bitaddie_4/xorg_0/m1_102_n17# 1bitaddie_4/Ai vdd 1bitaddie_4/xorg_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1242 1bitaddie_4/xorg_1/A 1bitaddie_4/xorg_0/inverter_1/out 1bitaddie_4/xorg_0/m1_102_n17# 1bitaddie_4/xorg_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 1bitaddie_4/xorg_1/inverter_0/out 1bitaddie_4/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1244 1bitaddie_4/xorg_1/inverter_0/out 1bitaddie_4/xorg_1/A vdd 1bitaddie_4/xorg_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1245 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/inverter_1/out gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1246 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/inverter_1/out vdd 1bitaddie_4/xorg_1/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1247 1bitaddie_4/sum 1bitaddie_4/inverter_1/out 1bitaddie_4/xorg_1/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1248 1bitaddie_4/xorg_1/m1_26_n95# 1bitaddie_4/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 1bitaddie_4/sum 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/xorg_1/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1250 1bitaddie_4/xorg_1/m1_102_n91# 1bitaddie_4/xorg_1/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 1bitaddie_4/xorg_1/m1_25_n11# 1bitaddie_4/xorg_1/inverter_0/out vdd 1bitaddie_4/xorg_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1252 1bitaddie_4/sum 1bitaddie_4/inverter_1/out 1bitaddie_4/xorg_1/m1_25_n11# 1bitaddie_4/xorg_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1253 1bitaddie_4/xorg_1/m1_102_n17# 1bitaddie_4/xorg_1/A vdd 1bitaddie_4/xorg_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1254 1bitaddie_4/sum 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/xorg_1/m1_102_n17# 1bitaddie_4/xorg_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 1bitaddie_4/Bi 1bitaddie_4/ff_0/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1256 1bitaddie_4/Bi 1bitaddie_4/ff_0/inverter_0/in vdd 1bitaddie_4/ff_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1257 1bitaddie_4/ff_0/m1_25_n37# B4 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1258 1bitaddie_4/ff_0/m1_63_0# 1bitaddie_4/ff_0/m1_25_n37# 1bitaddie_4/ff_0/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1259 1bitaddie_4/ff_0/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 1bitaddie_4/ff_0/inverter_0/in 1bitaddie_4/clk 1bitaddie_4/ff_0/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1261 1bitaddie_4/ff_0/m1_106_n52# 1bitaddie_4/ff_0/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1262 1bitaddie_4/ff_0/m1_19_n10# B4 vdd 1bitaddie_4/ff_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1263 1bitaddie_4/ff_0/m1_25_n37# 1bitaddie_4/clk 1bitaddie_4/ff_0/m1_19_n10# 1bitaddie_4/ff_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1264 1bitaddie_4/ff_0/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_4/ff_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1265 1bitaddie_4/ff_0/inverter_0/in 1bitaddie_4/ff_0/m1_63_0# vdd 1bitaddie_4/ff_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1266 1bitaddie_4/Ai 1bitaddie_4/ff_1/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1267 1bitaddie_4/Ai 1bitaddie_4/ff_1/inverter_0/in vdd 1bitaddie_4/ff_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1268 1bitaddie_4/ff_1/m1_25_n37# A4 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1269 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/ff_1/m1_25_n37# 1bitaddie_4/ff_1/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1270 1bitaddie_4/ff_1/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 1bitaddie_4/ff_1/inverter_0/in 1bitaddie_4/clk 1bitaddie_4/ff_1/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1272 1bitaddie_4/ff_1/m1_106_n52# 1bitaddie_4/ff_1/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 1bitaddie_4/ff_1/m1_19_n10# A4 vdd 1bitaddie_4/ff_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1274 1bitaddie_4/ff_1/m1_25_n37# 1bitaddie_4/clk 1bitaddie_4/ff_1/m1_19_n10# 1bitaddie_4/ff_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1275 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_4/ff_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1276 1bitaddie_4/ff_1/inverter_0/in 1bitaddie_4/ff_1/m1_63_0# vdd 1bitaddie_4/ff_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1277 s4 1bitaddie_4/ff_2/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1278 s4 1bitaddie_4/ff_2/inverter_0/in vdd 1bitaddie_4/ff_2/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1279 1bitaddie_4/ff_2/m1_25_n37# 1bitaddie_4/sum gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1280 1bitaddie_4/ff_2/m1_63_0# 1bitaddie_4/ff_2/m1_25_n37# 1bitaddie_4/ff_2/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1281 1bitaddie_4/ff_2/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1282 1bitaddie_4/ff_2/inverter_0/in 1bitaddie_4/clk 1bitaddie_4/ff_2/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1283 1bitaddie_4/ff_2/m1_106_n52# 1bitaddie_4/ff_2/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1284 1bitaddie_4/ff_2/m1_19_n10# 1bitaddie_4/sum vdd 1bitaddie_4/ff_2/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1285 1bitaddie_4/ff_2/m1_25_n37# 1bitaddie_4/clk 1bitaddie_4/ff_2/m1_19_n10# 1bitaddie_4/ff_2/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1286 1bitaddie_4/ff_2/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_4/ff_2/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1287 1bitaddie_4/ff_2/inverter_0/in 1bitaddie_4/ff_2/m1_63_0# vdd 1bitaddie_4/ff_2/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1288 inverter_0/in ff_0/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1289 inverter_0/in ff_0/inverter_0/in vdd ff_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1290 ff_0/m1_25_n37# C0 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1291 ff_0/m1_63_0# ff_0/m1_25_n37# ff_0/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1292 ff_0/m1_58_n52# m1_611_197# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1293 ff_0/inverter_0/in m1_560_235# ff_0/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1294 ff_0/m1_106_n52# ff_0/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 ff_0/m1_19_n10# C0 vdd ff_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1296 ff_0/m1_25_n37# m1_641_206# ff_0/m1_19_n10# ff_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1297 ff_0/m1_63_0# m1_608_244# vdd ff_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1298 ff_0/inverter_0/in ff_0/m1_63_0# vdd ff_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1299 Cout ff_1/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1300 Cout ff_1/inverter_0/in vdd ff_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1301 ff_1/m1_25_n37# inverter_1/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1302 ff_1/m1_63_0# ff_1/m1_25_n37# ff_1/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1303 ff_1/m1_58_n52# ff_1/nmos_2/a_0_n10# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 ff_1/inverter_0/in ff_1/nmos_3/a_0_n10# ff_1/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1305 ff_1/m1_106_n52# ff_1/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1306 ff_1/m1_19_n10# inverter_1/in vdd ff_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1307 ff_1/m1_25_n37# ff_1/pmos_1/a_0_n10# ff_1/m1_19_n10# ff_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1308 ff_1/m1_63_0# ff_1/pmos_2/a_0_n10# vdd ff_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1309 ff_1/inverter_0/in ff_1/m1_63_0# vdd ff_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1310 1bitaddie_0/inverter_0/in 1bitaddie_0/Bi 1bitaddie_0/nandg_0/m1_26_n48# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1311 1bitaddie_0/nandg_0/m1_26_n48# 1bitaddie_0/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1312 1bitaddie_0/inverter_0/in 1bitaddie_0/Bi vdd 1bitaddie_0/nandg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1313 1bitaddie_0/inverter_0/in 1bitaddie_0/Ai vdd 1bitaddie_0/nandg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1314 1bitaddie_0/inverter_0/out 1bitaddie_0/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1315 1bitaddie_0/inverter_0/out 1bitaddie_0/inverter_0/in vdd 1bitaddie_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1316 1bitaddie_0/inverter_1/out inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1317 1bitaddie_0/inverter_1/out inverter_0/out vdd 1bitaddie_0/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1318 1bitaddie_0/manch_0/clk 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1319 1bitaddie_0/manch_0/clk 1bitaddie_4/clk vdd 1bitaddie_0/inverter_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1320 1bitaddie_1/Cin 1bitaddie_0/inverter_0/out 1bitaddie_0/manch_0/m1_24_n50# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1321 1bitaddie_0/manch_0/m1_24_n50# 1bitaddie_0/manch_0/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 1bitaddie_1/Cin 1bitaddie_0/xorg_1/A inverter_0/out Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1323 1bitaddie_1/Cin 1bitaddie_0/manch_0/clk vdd 1bitaddie_0/manch_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1324 1bitaddie_0/xorg_0/inverter_0/out 1bitaddie_0/Ai gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1325 1bitaddie_0/xorg_0/inverter_0/out 1bitaddie_0/Ai vdd 1bitaddie_0/xorg_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1326 1bitaddie_0/xorg_0/inverter_1/out 1bitaddie_0/Bi gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1327 1bitaddie_0/xorg_0/inverter_1/out 1bitaddie_0/Bi vdd 1bitaddie_0/xorg_0/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1328 1bitaddie_0/xorg_1/A 1bitaddie_0/Bi 1bitaddie_0/xorg_0/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1329 1bitaddie_0/xorg_0/m1_26_n95# 1bitaddie_0/Ai gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1330 1bitaddie_0/xorg_1/A 1bitaddie_0/xorg_0/inverter_1/out 1bitaddie_0/xorg_0/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1331 1bitaddie_0/xorg_0/m1_102_n91# 1bitaddie_0/xorg_0/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1332 1bitaddie_0/xorg_0/m1_25_n11# 1bitaddie_0/xorg_0/inverter_0/out vdd 1bitaddie_0/xorg_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1333 1bitaddie_0/xorg_1/A 1bitaddie_0/Bi 1bitaddie_0/xorg_0/m1_25_n11# 1bitaddie_0/xorg_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1334 1bitaddie_0/xorg_0/m1_102_n17# 1bitaddie_0/Ai vdd 1bitaddie_0/xorg_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1335 1bitaddie_0/xorg_1/A 1bitaddie_0/xorg_0/inverter_1/out 1bitaddie_0/xorg_0/m1_102_n17# 1bitaddie_0/xorg_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 1bitaddie_0/xorg_1/inverter_0/out 1bitaddie_0/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1337 1bitaddie_0/xorg_1/inverter_0/out 1bitaddie_0/xorg_1/A vdd 1bitaddie_0/xorg_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1338 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/inverter_1/out gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1339 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/inverter_1/out vdd 1bitaddie_0/xorg_1/inverter_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1340 1bitaddie_0/sum 1bitaddie_0/inverter_1/out 1bitaddie_0/xorg_1/m1_26_n95# Gnd nfet w=4 l=2
+  ad=40 pd=36 as=40 ps=36
M1341 1bitaddie_0/xorg_1/m1_26_n95# 1bitaddie_0/xorg_1/A gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1342 1bitaddie_0/sum 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/xorg_1/m1_102_n91# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=40 ps=36
M1343 1bitaddie_0/xorg_1/m1_102_n91# 1bitaddie_0/xorg_1/inverter_0/out gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1344 1bitaddie_0/xorg_1/m1_25_n11# 1bitaddie_0/xorg_1/inverter_0/out vdd 1bitaddie_0/xorg_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1345 1bitaddie_0/sum 1bitaddie_0/inverter_1/out 1bitaddie_0/xorg_1/m1_25_n11# 1bitaddie_0/xorg_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1346 1bitaddie_0/xorg_1/m1_102_n17# 1bitaddie_0/xorg_1/A vdd 1bitaddie_0/xorg_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1347 1bitaddie_0/sum 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/xorg_1/m1_102_n17# 1bitaddie_0/xorg_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1348 1bitaddie_0/Bi 1bitaddie_0/ff_0/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1349 1bitaddie_0/Bi 1bitaddie_0/ff_0/inverter_0/in vdd 1bitaddie_0/ff_0/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1350 1bitaddie_0/ff_0/m1_25_n37# B0 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1351 1bitaddie_0/ff_0/m1_63_0# 1bitaddie_0/ff_0/m1_25_n37# 1bitaddie_0/ff_0/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1352 1bitaddie_0/ff_0/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1353 1bitaddie_0/ff_0/inverter_0/in 1bitaddie_4/clk 1bitaddie_0/ff_0/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1354 1bitaddie_0/ff_0/m1_106_n52# 1bitaddie_0/ff_0/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 1bitaddie_0/ff_0/m1_19_n10# B0 vdd 1bitaddie_0/ff_0/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1356 1bitaddie_0/ff_0/m1_25_n37# 1bitaddie_4/clk 1bitaddie_0/ff_0/m1_19_n10# 1bitaddie_0/ff_0/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1357 1bitaddie_0/ff_0/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_0/ff_0/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1358 1bitaddie_0/ff_0/inverter_0/in 1bitaddie_0/ff_0/m1_63_0# vdd 1bitaddie_0/ff_0/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1359 1bitaddie_0/Ai 1bitaddie_0/ff_1/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1360 1bitaddie_0/Ai 1bitaddie_0/ff_1/inverter_0/in vdd 1bitaddie_0/ff_1/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1361 1bitaddie_0/ff_1/m1_25_n37# A0 gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1362 1bitaddie_0/ff_1/m1_63_0# 1bitaddie_0/ff_1/m1_25_n37# 1bitaddie_0/ff_1/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1363 1bitaddie_0/ff_1/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1364 1bitaddie_0/ff_1/inverter_0/in 1bitaddie_4/clk 1bitaddie_0/ff_1/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1365 1bitaddie_0/ff_1/m1_106_n52# 1bitaddie_0/ff_1/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1366 1bitaddie_0/ff_1/m1_19_n10# A0 vdd 1bitaddie_0/ff_1/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1367 1bitaddie_0/ff_1/m1_25_n37# 1bitaddie_4/clk 1bitaddie_0/ff_1/m1_19_n10# 1bitaddie_0/ff_1/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1368 1bitaddie_0/ff_1/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_0/ff_1/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1369 1bitaddie_0/ff_1/inverter_0/in 1bitaddie_0/ff_1/m1_63_0# vdd 1bitaddie_0/ff_1/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1370 s0 1bitaddie_0/ff_2/inverter_0/in gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1371 s0 1bitaddie_0/ff_2/inverter_0/in vdd 1bitaddie_0/ff_2/inverter_0/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1372 1bitaddie_0/ff_2/m1_25_n37# 1bitaddie_0/sum gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1373 1bitaddie_0/ff_2/m1_63_0# 1bitaddie_0/ff_2/m1_25_n37# 1bitaddie_0/ff_2/m1_58_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1374 1bitaddie_0/ff_2/m1_58_n52# 1bitaddie_4/clk gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 1bitaddie_0/ff_2/inverter_0/in 1bitaddie_4/clk 1bitaddie_0/ff_2/m1_106_n52# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=40 ps=36
M1376 1bitaddie_0/ff_2/m1_106_n52# 1bitaddie_0/ff_2/m1_63_0# gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1377 1bitaddie_0/ff_2/m1_19_n10# 1bitaddie_0/sum vdd 1bitaddie_0/ff_2/pmos_0/w_n8_n5# pfet w=8 l=2
+  ad=80 pd=52 as=0 ps=0
M1378 1bitaddie_0/ff_2/m1_25_n37# 1bitaddie_4/clk 1bitaddie_0/ff_2/m1_19_n10# 1bitaddie_0/ff_2/pmos_1/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1379 1bitaddie_0/ff_2/m1_63_0# 1bitaddie_4/clk vdd 1bitaddie_0/ff_2/pmos_2/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1380 1bitaddie_0/ff_2/inverter_0/in 1bitaddie_0/ff_2/m1_63_0# vdd 1bitaddie_0/ff_2/pmos_3/w_n8_n5# pfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
C0 1bitaddie_4/clk 1bitaddie_0/ff_0/pmos_1/w_n8_n5# 0.30fF
C1 1bitaddie_2/xorg_0/m1_25_n11# 1bitaddie_2/xorg_1/A 0.12fF
C2 ff_1/inverter_0/w_n8_n5# Cout 0.03fF
C3 1bitaddie_0/Ai gnd 0.27fF
C4 1bitaddie_0/manch_0/m1_24_n50# gnd 0.08fF
C5 ff_1/pmos_2/w_n8_n5# ff_1/pmos_2/a_0_n10# 0.07fF
C6 1bitaddie_3/ff_1/pmos_3/w_n8_n5# vdd 0.06fF
C7 gnd 1bitaddie_3/nandg_0/m1_26_n48# 0.08fF
C8 1bitaddie_4/clk 1bitaddie_1/ff_2/m1_63_0# 0.27fF
C9 1bitaddie_3/ff_1/m1_25_n37# 1bitaddie_4/clk 0.41fF
C10 1bitaddie_0/xorg_0/inverter_1/out gnd 0.08fF
C11 1bitaddie_1/xorg_0/m1_25_n11# 1bitaddie_1/xorg_1/A 0.12fF
C12 1bitaddie_4/ff_1/pmos_1/w_n8_n5# 1bitaddie_4/ff_1/m1_25_n37# 0.03fF
C13 inverter_0/in gnd 0.14fF
C14 B2 1bitaddie_2/ff_0/pmos_0/w_n8_n5# 0.07fF
C15 1bitaddie_0/ff_0/m1_19_n10# vdd 0.12fF
C16 1bitaddie_3/inverter_1/out gnd 0.14fF
C17 1bitaddie_1/ff_2/m1_106_n52# 1bitaddie_1/ff_2/m1_63_0# 0.05fF
C18 A0 1bitaddie_0/ff_1/m1_19_n10# 0.11fF
C19 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/clk 0.35fF
C20 1bitaddie_3/ff_2/inverter_0/in s3 0.05fF
C21 1bitaddie_0/manch_0/pmos_0/w_n8_n5# 1bitaddie_0/manch_0/clk 0.07fF
C22 inverter_1/in ff_1/pmos_1/a_0_n10# 0.05fF
C23 1bitaddie_4/Bi gnd 0.18fF
C24 1bitaddie_4/nandg_0/pmos_1/w_n8_n5# vdd 0.08fF
C25 gnd 1bitaddie_1/xorg_1/inverter_0/out 0.14fF
C26 1bitaddie_0/xorg_1/inverter_1/out gnd 0.08fF
C27 1bitaddie_2/xorg_1/inverter_0/w_n8_n5# 1bitaddie_2/xorg_1/inverter_0/out 0.03fF
C28 1bitaddie_1/ff_2/m1_58_n52# 1bitaddie_1/ff_2/m1_63_0# 0.08fF
C29 1bitaddie_2/sum 1bitaddie_2/ff_2/m1_25_n37# 0.05fF
C30 1bitaddie_3/xorg_1/inverter_0/out 1bitaddie_3/xorg_1/m1_25_n11# 0.05fF
C31 gnd 1bitaddie_1/xorg_1/m1_102_n91# 0.08fF
C32 1bitaddie_4/xorg_1/inverter_0/w_n8_n5# 1bitaddie_4/xorg_1/A 0.07fF
C33 1bitaddie_4/manch_0/clk 1bitaddie_4/clk 0.05fF
C34 1bitaddie_3/xorg_0/inverter_0/out 1bitaddie_3/xorg_1/A 0.06fF
C35 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/xorg_1/inverter_1/w_n8_n5# 0.03fF
C36 1bitaddie_0/xorg_0/inverter_0/out 1bitaddie_0/xorg_0/m1_25_n11# 0.05fF
C37 1bitaddie_4/nandg_0/m1_26_n48# gnd 0.08fF
C38 1bitaddie_2/xorg_1/A 1bitaddie_2/xorg_1/m1_102_n17# 0.20fF
C39 1bitaddie_1/Ai 1bitaddie_1/Bi 0.06fF
C40 gnd A1 0.05fF
C41 1bitaddie_2/inverter_0/out vdd 0.12fF
C42 1bitaddie_3/xorg_0/m1_25_n11# 1bitaddie_3/xorg_1/A 0.12fF
C43 1bitaddie_2/ff_2/pmos_3/w_n8_n5# vdd 0.06fF
C44 1bitaddie_4/xorg_1/pmos_3/w_n8_n5# 1bitaddie_4/xorg_1/m1_102_n17# 0.08fF
C45 1bitaddie_2/ff_2/m1_25_n37# 1bitaddie_4/clk 0.27fF
C46 1bitaddie_2/ff_0/m1_58_n52# 1bitaddie_4/clk 0.12fF
C47 gnd 1bitaddie_1/ff_0/m1_25_n37# 0.08fF
C48 1bitaddie_1/inverter_0/out 1bitaddie_1/manch_0/clk 0.03fF
C49 1bitaddie_0/xorg_1/m1_26_n95# gnd 0.08fF
C50 1bitaddie_4/ff_2/pmos_1/w_n8_n5# 1bitaddie_4/ff_2/m1_19_n10# 0.08fF
C51 1bitaddie_4/Cin 1bitaddie_4/clk 0.11fF
C52 inverter_1/out vdd 0.25fF
C53 1bitaddie_3/inverter_0/in 1bitaddie_3/nandg_0/pmos_1/w_n8_n5# 0.03fF
C54 1bitaddie_2/ff_0/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.30fF
C55 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/sum 0.22fF
C56 1bitaddie_4/clk 1bitaddie_0/ff_1/pmos_1/w_n8_n5# 0.31fF
C57 1bitaddie_4/Bi 1bitaddie_4/ff_0/inverter_0/w_n8_n5# 0.03fF
C58 B3 1bitaddie_3/ff_0/pmos_0/w_n8_n5# 0.07fF
C59 1bitaddie_2/Ai gnd 0.27fF
C60 1bitaddie_0/xorg_1/A gnd 0.48fF
C61 1bitaddie_2/manch_0/m1_24_n50# gnd 0.08fF
C62 1bitaddie_0/ff_2/inverter_0/in 1bitaddie_0/ff_2/inverter_0/w_n8_n5# 0.07fF
C63 1bitaddie_3/inverter_2/w_n8_n5# vdd 0.08fF
C64 1bitaddie_3/inverter_0/out vdd 0.12fF
C65 1bitaddie_3/ff_2/pmos_3/w_n8_n5# vdd 0.06fF
C66 ff_1/m1_63_0# vdd 0.12fF
C67 1bitaddie_3/ff_2/m1_25_n37# 1bitaddie_4/clk 0.27fF
C68 1bitaddie_3/ff_0/m1_58_n52# 1bitaddie_4/clk 0.12fF
C69 1bitaddie_3/xorg_1/inverter_0/w_n8_n5# 1bitaddie_3/xorg_1/inverter_0/out 0.03fF
C70 1bitaddie_2/xorg_0/inverter_1/out gnd 0.08fF
C71 1bitaddie_4/xorg_0/inverter_0/out gnd 0.14fF
C72 1bitaddie_3/sum 1bitaddie_3/ff_2/m1_25_n37# 0.05fF
C73 1bitaddie_2/ff_0/m1_19_n10# vdd 0.12fF
C74 1bitaddie_0/ff_1/m1_19_n10# vdd 0.12fF
C75 vdd 1bitaddie_1/xorg_1/inverter_1/out 0.12fF
C76 1bitaddie_3/ff_0/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.30fF
C77 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/xorg_1/inverter_1/w_n8_n5# 0.03fF
C78 1bitaddie_1/xorg_0/inverter_1/out 1bitaddie_1/xorg_0/m1_102_n91# 0.05fF
C79 1bitaddie_4/inverter_0/in 1bitaddie_4/nandg_0/pmos_1/w_n8_n5# 0.03fF
C80 1bitaddie_2/xorg_1/inverter_1/out gnd 0.08fF
C81 1bitaddie_1/manch_0/clk 1bitaddie_4/clk 0.05fF
C82 1bitaddie_4/nandg_0/pmos_0/w_n8_n5# vdd 0.08fF
C83 1bitaddie_3/xorg_1/A 1bitaddie_3/xorg_1/m1_102_n17# 0.20fF
C84 1bitaddie_3/Ai gnd 0.27fF
C85 1bitaddie_2/ff_0/m1_19_n10# 1bitaddie_2/ff_0/m1_25_n37# 0.12fF
C86 1bitaddie_4/inverter_1/out 1bitaddie_4/xorg_1/pmos_1/w_n8_n5# 0.07fF
C87 1bitaddie_3/manch_0/m1_24_n50# gnd 0.08fF
C88 1bitaddie_4/clk 1bitaddie_0/ff_1/inverter_0/in 0.05fF
C89 1bitaddie_4/sum 1bitaddie_4/xorg_1/m1_26_n95# 0.08fF
C90 1bitaddie_0/ff_1/m1_19_n10# 1bitaddie_0/ff_1/m1_25_n37# 0.12fF
C91 ff_0/pmos_2/w_n8_n5# vdd 0.08fF
C92 1bitaddie_4/ff_0/pmos_0/w_n8_n5# vdd 0.08fF
C93 1bitaddie_0/Ai 1bitaddie_0/ff_1/inverter_0/w_n8_n5# 0.03fF
C94 1bitaddie_3/xorg_0/inverter_1/out gnd 0.08fF
C95 1bitaddie_0/ff_1/inverter_0/in 1bitaddie_0/ff_1/pmos_3/w_n8_n5# 0.03fF
C96 Cout gnd 0.08fF
C97 1bitaddie_0/ff_0/pmos_1/w_n8_n5# 1bitaddie_0/ff_0/m1_19_n10# 0.08fF
C98 1bitaddie_0/ff_0/pmos_0/w_n8_n5# 1bitaddie_0/ff_0/m1_19_n10# 0.03fF
C99 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/xorg_1/pmos_3/w_n8_n5# 0.07fF
C100 1bitaddie_0/xorg_0/pmos_1/w_n8_n5# 1bitaddie_0/xorg_1/A 0.03fF
C101 1bitaddie_3/ff_0/m1_19_n10# vdd 0.12fF
C102 gnd 1bitaddie_1/xorg_0/m1_102_n91# 0.08fF
C103 A0 1bitaddie_0/ff_1/m1_25_n37# 0.05fF
C104 1bitaddie_1/Ai 1bitaddie_1/xorg_0/m1_25_n11# 0.14fF
C105 1bitaddie_3/xorg_1/inverter_1/out gnd 0.08fF
C106 1bitaddie_4/xorg_0/inverter_0/w_n8_n5# 1bitaddie_4/xorg_0/inverter_0/out 0.03fF
C107 1bitaddie_0/ff_0/m1_63_0# 1bitaddie_0/ff_0/pmos_2/w_n8_n5# 0.03fF
C108 1bitaddie_2/xorg_1/m1_26_n95# gnd 0.08fF
C109 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/ff_1/m1_25_n37# 0.05fF
C110 1bitaddie_0/nandg_0/pmos_0/w_n8_n5# 1bitaddie_0/Bi 0.07fF
C111 ff_1/pmos_0/w_n8_n5# vdd 0.08fF
C112 1bitaddie_2/ff_1/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.31fF
C113 1bitaddie_1/ff_2/m1_25_n37# gnd 0.08fF
C114 1bitaddie_4/clk 1bitaddie_0/ff_2/pmos_1/w_n8_n5# 0.07fF
C115 1bitaddie_2/xorg_1/A gnd 0.48fF
C116 1bitaddie_1/xorg_0/inverter_0/out gnd 0.14fF
C117 1bitaddie_4/Ai 1bitaddie_4/xorg_0/m1_26_n95# 0.05fF
C118 inverter_0/in ff_0/inverter_0/w_n8_n5# 0.03fF
C119 1bitaddie_4/xorg_0/inverter_1/w_n8_n5# 1bitaddie_4/Bi 0.07fF
C120 1bitaddie_3/ff_0/m1_19_n10# 1bitaddie_3/ff_0/m1_25_n37# 0.12fF
C121 1bitaddie_0/xorg_0/pmos_2/w_n8_n5# vdd 0.08fF
C122 1bitaddie_3/nandg_0/pmos_0/w_n8_n5# 1bitaddie_3/Bi 0.07fF
C123 1bitaddie_1/sum 1bitaddie_1/xorg_1/pmos_1/w_n8_n5# 0.03fF
C124 inverter_0/w_n8_n5# inverter_0/out 0.03fF
C125 1bitaddie_4/ff_0/m1_106_n52# gnd 0.08fF
C126 1bitaddie_3/xorg_1/m1_26_n95# gnd 0.08fF
C127 1bitaddie_4/ff_2/pmos_1/w_n8_n5# 1bitaddie_4/ff_2/m1_25_n37# 0.03fF
C128 A2 1bitaddie_2/ff_1/m1_19_n10# 0.11fF
C129 1bitaddie_2/ff_1/m1_19_n10# vdd 0.12fF
C130 1bitaddie_4/xorg_1/inverter_0/out vdd 0.12fF
C131 1bitaddie_2/manch_0/pmos_0/w_n8_n5# 1bitaddie_2/manch_0/clk 0.07fF
C132 1bitaddie_2/nandg_0/pmos_0/w_n8_n5# 1bitaddie_2/inverter_0/in 0.03fF
C133 vdd 1bitaddie_0/ff_2/m1_19_n10# 0.12fF
C134 vdd 1bitaddie_1/ff_0/m1_63_0# 0.12fF
C135 1bitaddie_3/ff_1/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.31fF
C136 1bitaddie_4/inverter_0/in 1bitaddie_4/nandg_0/pmos_0/w_n8_n5# 0.03fF
C137 1bitaddie_3/xorg_1/A gnd 0.48fF
C138 vdd 1bitaddie_1/ff_1/pmos_0/w_n8_n5# 0.08fF
C139 1bitaddie_1/xorg_1/inverter_0/out 1bitaddie_1/xorg_1/pmos_0/w_n8_n5# 0.07fF
C140 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/inverter_1/out 0.05fF
C141 1bitaddie_2/ff_1/inverter_0/in 1bitaddie_4/clk 0.05fF
C142 gnd B1 0.05fF
C143 1bitaddie_1/Ai 1bitaddie_1/ff_1/inverter_0/in 0.05fF
C144 ff_0/m1_106_n52# ff_0/m1_63_0# 0.05fF
C145 1bitaddie_4/ff_2/m1_63_0# 1bitaddie_4/ff_2/pmos_2/w_n8_n5# 0.03fF
C146 vdd 1bitaddie_1/xorg_1/inverter_0/w_n8_n5# 0.08fF
C147 1bitaddie_2/xorg_0/inverter_0/out 1bitaddie_2/xorg_0/m1_25_n11# 0.05fF
C148 1bitaddie_1/Cin 1bitaddie_1/inverter_1/w_n8_n5# 0.07fF
C149 1bitaddie_3/ff_1/m1_19_n10# vdd 0.12fF
C150 gnd 1bitaddie_1/ff_1/m1_63_0# 0.05fF
C151 1bitaddie_4/clk 1bitaddie_0/ff_1/m1_63_0# 0.35fF
C152 1bitaddie_0/Bi gnd 0.18fF
C153 1bitaddie_3/ff_1/inverter_0/in 1bitaddie_4/clk 0.05fF
C154 1bitaddie_0/ff_1/m1_63_0# 1bitaddie_0/ff_1/pmos_3/w_n8_n5# 0.07fF
C155 1bitaddie_4/manch_0/clk inverter_1/out 0.16fF
C156 1bitaddie_1/xorg_1/pmos_2/w_n8_n5# 1bitaddie_1/xorg_1/m1_102_n17# 0.03fF
C157 1bitaddie_1/Bi A1 0.03fF
C158 1bitaddie_0/ff_0/m1_58_n52# 1bitaddie_0/ff_0/m1_25_n37# 0.08fF
C159 1bitaddie_4/ff_1/inverter_0/in vdd 0.12fF
C160 1bitaddie_4/Bi 1bitaddie_4/ff_0/inverter_0/in 0.05fF
C161 1bitaddie_2/manch_0/pmos_0/w_n8_n5# 1bitaddie_3/Cin 0.03fF
C162 1bitaddie_2/ff_2/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.07fF
C163 1bitaddie_0/ff_0/pmos_1/w_n8_n5# 1bitaddie_0/ff_0/m1_25_n37# 0.03fF
C164 1bitaddie_0/xorg_0/inverter_0/w_n8_n5# 1bitaddie_0/Ai 0.07fF
C165 1bitaddie_4/clk 1bitaddie_0/manch_0/clk 0.05fF
C166 1bitaddie_4/ff_1/m1_106_n52# gnd 0.08fF
C167 A3 1bitaddie_3/ff_1/m1_19_n10# 0.11fF
C168 gnd s1 0.08fF
C169 1bitaddie_3/manch_0/pmos_0/w_n8_n5# 1bitaddie_3/manch_0/clk 0.07fF
C170 1bitaddie_4/inverter_0/out 1bitaddie_4/manch_0/m1_24_n50# 0.05fF
C171 1bitaddie_2/ff_2/inverter_0/in 1bitaddie_2/ff_2/inverter_0/w_n8_n5# 0.07fF
C172 1bitaddie_4/xorg_0/pmos_2/w_n8_n5# 1bitaddie_4/xorg_0/m1_102_n17# 0.03fF
C173 1bitaddie_4/xorg_0/m1_26_n95# 1bitaddie_4/xorg_1/A 0.08fF
C174 1bitaddie_4/clk 1bitaddie_1/ff_0/m1_58_n52# 0.12fF
C175 inverter_1/out 1bitaddie_4/Cin 0.14fF
C176 1bitaddie_1/inverter_0/out 1bitaddie_1/xorg_1/A 0.06fF
C177 1bitaddie_2/xorg_0/pmos_2/w_n8_n5# vdd 0.08fF
C178 1bitaddie_4/ff_1/m1_58_n52# gnd 0.08fF
C179 1bitaddie_4/inverter_1/out 1bitaddie_4/clk 0.06fF
C180 vdd 1bitaddie_1/ff_2/inverter_0/in 0.12fF
C181 1bitaddie_1/xorg_1/pmos_0/w_n8_n5# 1bitaddie_1/xorg_1/m1_25_n11# 0.03fF
C182 1bitaddie_0/xorg_1/m1_102_n91# 1bitaddie_0/sum 0.08fF
C183 1bitaddie_4/ff_0/m1_63_0# gnd 0.05fF
C184 1bitaddie_0/Bi 1bitaddie_0/xorg_0/pmos_1/w_n8_n5# 0.07fF
C185 1bitaddie_2/ff_2/m1_19_n10# vdd 0.12fF
C186 1bitaddie_3/inverter_0/out 1bitaddie_4/Cin 0.19fF
C187 1bitaddie_3/xorg_0/inverter_0/out 1bitaddie_3/xorg_0/m1_25_n11# 0.05fF
C188 1bitaddie_4/xorg_1/pmos_0/w_n8_n5# 1bitaddie_4/xorg_1/m1_25_n11# 0.03fF
C189 1bitaddie_3/ff_2/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.07fF
C190 1bitaddie_1/xorg_0/inverter_0/w_n8_n5# 1bitaddie_1/xorg_0/inverter_0/out 0.03fF
C191 1bitaddie_4/ff_2/inverter_0/in 1bitaddie_4/ff_2/m1_106_n52# 0.08fF
C192 vdd 1bitaddie_1/ff_2/pmos_0/w_n8_n5# 0.08fF
C193 1bitaddie_1/nandg_0/pmos_1/w_n8_n5# 1bitaddie_1/Ai 0.07fF
C194 1bitaddie_2/ff_1/m1_19_n10# 1bitaddie_2/ff_1/m1_25_n37# 0.12fF
C195 ff_1/nmos_2/a_0_n10# ff_1/m1_58_n52# 0.05fF
C196 1bitaddie_2/Ai 1bitaddie_2/ff_1/inverter_0/w_n8_n5# 0.03fF
C197 1bitaddie_1/xorg_1/m1_26_n95# 1bitaddie_1/xorg_1/A 0.05fF
C198 1bitaddie_4/clk 1bitaddie_1/ff_0/inverter_0/in 0.22fF
C199 1bitaddie_0/ff_2/m1_19_n10# 1bitaddie_0/ff_2/m1_25_n37# 0.12fF
C200 1bitaddie_0/ff_0/m1_106_n52# 1bitaddie_0/ff_0/m1_63_0# 0.05fF
C201 1bitaddie_4/inverter_0/in vdd 0.25fF
C202 1bitaddie_3/xorg_0/pmos_2/w_n8_n5# vdd 0.08fF
C203 1bitaddie_2/ff_1/inverter_0/in 1bitaddie_2/ff_1/pmos_3/w_n8_n5# 0.03fF
C204 1bitaddie_2/ff_0/pmos_1/w_n8_n5# 1bitaddie_2/ff_0/m1_19_n10# 0.08fF
C205 1bitaddie_2/ff_0/pmos_0/w_n8_n5# 1bitaddie_2/ff_0/m1_19_n10# 0.03fF
C206 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/xorg_1/pmos_3/w_n8_n5# 0.07fF
C207 1bitaddie_2/xorg_0/pmos_1/w_n8_n5# 1bitaddie_2/xorg_1/A 0.03fF
C208 vdd 1bitaddie_1/inverter_1/out 0.18fF
C209 1bitaddie_0/xorg_0/inverter_0/out gnd 0.14fF
C210 1bitaddie_0/ff_1/pmos_1/w_n8_n5# 1bitaddie_0/ff_1/m1_19_n10# 0.08fF
C211 1bitaddie_3/ff_2/m1_19_n10# vdd 0.12fF
C212 1bitaddie_4/clk 1bitaddie_1/xorg_1/A 0.06fF
C213 A2 1bitaddie_2/ff_1/m1_25_n37# 0.05fF
C214 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_4/clk 0.35fF
C215 1bitaddie_2/Bi gnd 0.18fF
C216 1bitaddie_1/inverter_0/out 1bitaddie_2/Cin 0.19fF
C217 gnd 1bitaddie_1/Cin 0.10fF
C218 1bitaddie_2/ff_0/m1_63_0# 1bitaddie_2/ff_0/pmos_2/w_n8_n5# 0.03fF
C219 1bitaddie_3/ff_2/inverter_0/in 1bitaddie_3/ff_2/inverter_0/w_n8_n5# 0.07fF
C220 1bitaddie_1/xorg_0/pmos_1/w_n8_n5# 1bitaddie_1/xorg_1/A 0.03fF
C221 vdd 1bitaddie_1/ff_0/inverter_0/w_n8_n5# 0.08fF
C222 1bitaddie_0/ff_0/pmos_0/w_n8_n5# vdd 0.08fF
C223 1bitaddie_2/manch_0/clk 1bitaddie_4/clk 0.05fF
C224 ff_1/pmos_1/a_0_n10# ff_1/m1_25_n37# 0.05fF
C225 1bitaddie_4/inverter_0/out 1bitaddie_4/xorg_1/A 0.06fF
C226 1bitaddie_4/ff_2/m1_106_n52# gnd 0.08fF
C227 1bitaddie_4/ff_2/m1_63_0# 1bitaddie_4/ff_2/m1_106_n52# 0.05fF
C228 s4 vdd 0.12fF
C229 vdd 1bitaddie_1/ff_2/m1_63_0# 0.12fF
C230 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_4/clk 0.35fF
C231 1bitaddie_3/Bi gnd 0.18fF
C232 1bitaddie_0/inverter_0/out 1bitaddie_0/manch_0/clk 0.03fF
C233 inverter_1/in inverter_1/out 0.05fF
C234 gnd 1bitaddie_1/sum 0.35fF
C235 ff_1/m1_63_0# ff_1/pmos_3/w_n8_n5# 0.07fF
C236 1bitaddie_4/ff_1/m1_63_0# vdd 0.12fF
C237 1bitaddie_3/ff_1/m1_19_n10# 1bitaddie_3/ff_1/m1_25_n37# 0.12fF
C238 1bitaddie_4/ff_2/m1_58_n52# gnd 0.08fF
C239 1bitaddie_4/ff_2/m1_63_0# 1bitaddie_4/ff_2/m1_58_n52# 0.08fF
C240 1bitaddie_3/Ai 1bitaddie_3/ff_1/inverter_0/w_n8_n5# 0.03fF
C241 1bitaddie_2/Cin 1bitaddie_4/clk 0.11fF
C242 1bitaddie_0/inverter_1/out 1bitaddie_0/sum 0.20fF
C243 1bitaddie_4/inverter_0/w_n8_n5# 1bitaddie_4/inverter_0/out 0.03fF
C244 1bitaddie_3/ff_1/inverter_0/in 1bitaddie_3/ff_1/pmos_3/w_n8_n5# 0.03fF
C245 1bitaddie_1/nandg_0/pmos_0/w_n8_n5# 1bitaddie_1/Bi 0.07fF
C246 1bitaddie_0/xorg_0/pmos_1/w_n8_n5# 1bitaddie_0/xorg_0/m1_25_n11# 0.08fF
C247 1bitaddie_3/ff_0/pmos_1/w_n8_n5# 1bitaddie_3/ff_0/m1_19_n10# 0.08fF
C248 1bitaddie_3/ff_0/pmos_0/w_n8_n5# 1bitaddie_3/ff_0/m1_19_n10# 0.03fF
C249 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/xorg_1/pmos_3/w_n8_n5# 0.07fF
C250 1bitaddie_3/xorg_0/pmos_1/w_n8_n5# 1bitaddie_3/xorg_1/A 0.03fF
C251 1bitaddie_3/manch_0/clk 1bitaddie_4/clk 0.05fF
C252 1bitaddie_0/inverter_0/out inverter_0/out 0.02fF
C253 1bitaddie_0/xorg_0/inverter_1/w_n8_n5# 1bitaddie_0/xorg_0/inverter_1/out 0.03fF
C254 ff_1/m1_58_n52# ff_1/m1_25_n37# 0.08fF
C255 A3 1bitaddie_3/ff_1/m1_25_n37# 0.05fF
C256 1bitaddie_4/manch_0/clk vdd 0.12fF
C257 ff_0/pmos_3/w_n8_n5# vdd 0.06fF
C258 1bitaddie_3/ff_0/m1_63_0# 1bitaddie_3/ff_0/pmos_2/w_n8_n5# 0.03fF
C259 1bitaddie_3/nandg_0/pmos_1/w_n8_n5# vdd 0.08fF
C260 1bitaddie_4/clk 1bitaddie_1/ff_1/m1_19_n10# 0.09fF
C261 gnd 1bitaddie_1/inverter_0/in 0.05fF
C262 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/ff_1/inverter_0/in 0.05fF
C263 1bitaddie_1/ff_1/inverter_0/w_n8_n5# 1bitaddie_1/Ai 0.03fF
C264 1bitaddie_0/ff_0/m1_106_n52# gnd 0.08fF
C265 1bitaddie_3/Cin 1bitaddie_4/clk 0.11fF
C266 1bitaddie_2/xorg_0/inverter_0/out gnd 0.14fF
C267 1bitaddie_1/xorg_1/A 1bitaddie_1/xorg_1/pmos_2/w_n8_n5# 0.07fF
C268 1bitaddie_1/inverter_0/out 1bitaddie_1/manch_0/m1_24_n50# 0.05fF
C269 1bitaddie_0/inverter_1/w_n8_n5# vdd 0.08fF
C270 ff_0/inverter_0/in ff_0/m1_63_0# 0.05fF
C271 1bitaddie_1/xorg_0/pmos_3/w_n8_n5# 1bitaddie_1/xorg_0/m1_102_n17# 0.08fF
C272 1bitaddie_0/xorg_1/inverter_0/out vdd 0.12fF
C273 1bitaddie_1/ff_2/inverter_0/in 1bitaddie_1/ff_2/m1_63_0# 0.05fF
C274 1bitaddie_4/Cin vdd 0.12fF
C275 1bitaddie_0/xorg_1/A 1bitaddie_0/xorg_1/m1_25_n11# 0.14fF
C276 1bitaddie_4/Bi 1bitaddie_4/xorg_0/m1_26_n95# 0.05fF
C277 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_2/ff_1/pmos_3/w_n8_n5# 0.07fF
C278 1bitaddie_4/ff_0/inverter_0/in 1bitaddie_4/ff_0/m1_106_n52# 0.08fF
C279 1bitaddie_2/ff_0/m1_58_n52# 1bitaddie_2/ff_0/m1_25_n37# 0.08fF
C280 1bitaddie_0/nandg_0/m1_26_n48# 1bitaddie_0/inverter_0/in 0.08fF
C281 1bitaddie_2/ff_0/pmos_0/w_n8_n5# vdd 0.08fF
C282 1bitaddie_2/ff_0/pmos_1/w_n8_n5# 1bitaddie_2/ff_0/m1_25_n37# 0.03fF
C283 1bitaddie_2/xorg_0/inverter_0/w_n8_n5# 1bitaddie_2/Ai 0.07fF
C284 1bitaddie_4/sum 1bitaddie_4/xorg_1/m1_102_n17# 0.12fF
C285 1bitaddie_3/xorg_0/inverter_0/out gnd 0.14fF
C286 1bitaddie_0/ff_1/pmos_1/w_n8_n5# 1bitaddie_0/ff_1/m1_25_n37# 0.03fF
C287 ff_0/m1_19_n10# vdd 0.12fF
C288 C0 gnd 0.05fF
C289 ff_0/m1_58_n52# m1_611_197# 0.05fF
C290 inverter_1/in ff_1/pmos_0/w_n8_n5# 0.07fF
C291 1bitaddie_3/ff_0/pmos_0/w_n8_n5# vdd 0.08fF
C292 1bitaddie_2/xorg_1/m1_102_n91# 1bitaddie_2/sum 0.08fF
C293 1bitaddie_2/Bi 1bitaddie_2/xorg_0/pmos_1/w_n8_n5# 0.07fF
C294 1bitaddie_1/xorg_0/inverter_0/out 1bitaddie_1/xorg_0/m1_25_n11# 0.05fF
C295 1bitaddie_1/manch_0/clk vdd 0.12fF
C296 s1 1bitaddie_1/ff_2/inverter_0/w_n8_n5# 0.03fF
C297 1bitaddie_0/ff_1/inverter_0/in vdd 0.12fF
C298 1bitaddie_4/xorg_1/A 1bitaddie_4/clk 0.06fF
C299 1bitaddie_0/xorg_1/inverter_0/w_n8_n5# 1bitaddie_0/xorg_1/A 0.07fF
C300 1bitaddie_0/ff_1/m1_106_n52# gnd 0.08fF
C301 ff_1/m1_63_0# ff_1/pmos_2/a_0_n10# 0.05fF
C302 1bitaddie_4/Ai 1bitaddie_4/xorg_0/pmos_2/w_n8_n5# 0.07fF
C303 1bitaddie_2/ff_2/m1_19_n10# 1bitaddie_2/ff_2/m1_25_n37# 0.12fF
C304 1bitaddie_2/ff_0/m1_106_n52# 1bitaddie_2/ff_0/m1_63_0# 0.05fF
C305 ff_1/pmos_3/w_n8_n5# vdd 0.06fF
C306 ff_0/pmos_1/w_n8_n5# ff_0/m1_19_n10# 0.08fF
C307 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_3/ff_1/pmos_3/w_n8_n5# 0.07fF
C308 1bitaddie_3/ff_0/m1_58_n52# 1bitaddie_3/ff_0/m1_25_n37# 0.08fF
C309 1bitaddie_0/ff_1/m1_58_n52# gnd 0.08fF
C310 1bitaddie_4/clk 1bitaddie_0/inverter_1/out 0.06fF
C311 1bitaddie_0/xorg_1/pmos_3/w_n8_n5# 1bitaddie_0/xorg_1/m1_102_n17# 0.08fF
C312 1bitaddie_2/ff_1/pmos_1/w_n8_n5# 1bitaddie_2/ff_1/m1_19_n10# 0.08fF
C313 1bitaddie_2/ff_0/m1_106_n52# gnd 0.08fF
C314 1bitaddie_0/ff_2/pmos_1/w_n8_n5# 1bitaddie_0/ff_2/m1_19_n10# 0.08fF
C315 1bitaddie_0/ff_0/m1_63_0# gnd 0.05fF
C316 1bitaddie_2/xorg_1/inverter_0/out vdd 0.12fF
C317 1bitaddie_3/ff_0/pmos_1/w_n8_n5# 1bitaddie_3/ff_0/m1_25_n37# 0.03fF
C318 1bitaddie_3/xorg_0/inverter_0/w_n8_n5# 1bitaddie_3/Ai 0.07fF
C319 vdd 1bitaddie_1/xorg_1/m1_102_n17# 0.12fF
C320 1bitaddie_2/nandg_0/pmos_1/w_n8_n5# 1bitaddie_2/inverter_0/in 0.03fF
C321 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/sum 0.22fF
C322 1bitaddie_0/Bi 1bitaddie_0/ff_0/inverter_0/w_n8_n5# 0.03fF
C323 1bitaddie_4/xorg_1/m1_102_n91# 1bitaddie_4/xorg_1/inverter_0/out 0.05fF
C324 1bitaddie_4/xorg_0/m1_102_n17# vdd 0.12fF
C325 1bitaddie_4/ff_0/inverter_0/in 1bitaddie_4/ff_0/m1_63_0# 0.05fF
C326 1bitaddie_4/xorg_0/pmos_0/w_n8_n5# vdd 0.08fF
C327 inverter_0/in inverter_0/w_n8_n5# 0.07fF
C328 inverter_0/in ff_0/inverter_0/in 0.05fF
C329 vdd 1bitaddie_1/ff_1/pmos_3/w_n8_n5# 0.06fF
C330 1bitaddie_1/inverter_0/w_n8_n5# 1bitaddie_1/inverter_0/in 0.07fF
C331 1bitaddie_4/clk 1bitaddie_1/ff_1/m1_25_n37# 0.41fF
C332 1bitaddie_3/ff_0/m1_106_n52# gnd 0.08fF
C333 1bitaddie_3/xorg_1/m1_102_n91# 1bitaddie_3/sum 0.08fF
C334 1bitaddie_3/Bi 1bitaddie_3/xorg_0/pmos_1/w_n8_n5# 0.07fF
C335 ff_0/m1_58_n52# ff_0/m1_25_n37# 0.08fF
C336 1bitaddie_3/xorg_1/inverter_0/out vdd 0.12fF
C337 1bitaddie_4/nandg_0/pmos_1/w_n8_n5# 1bitaddie_4/Ai 0.07fF
C338 1bitaddie_2/inverter_0/out 1bitaddie_2/manch_0/clk 0.03fF
C339 1bitaddie_4/clk 1bitaddie_1/ff_0/m1_19_n10# 0.09fF
C340 1bitaddie_4/ff_2/inverter_0/in 1bitaddie_4/ff_2/m1_63_0# 0.05fF
C341 1bitaddie_4/ff_2/inverter_0/in gnd 0.05fF
C342 1bitaddie_1/Bi 1bitaddie_1/xorg_0/m1_102_n17# 0.05fF
C343 ff_1/pmos_1/w_n8_n5# ff_1/pmos_1/a_0_n10# 0.07fF
C344 1bitaddie_3/ff_2/m1_19_n10# 1bitaddie_3/ff_2/m1_25_n37# 0.12fF
C345 1bitaddie_0/inverter_1/out 1bitaddie_0/xorg_1/pmos_1/w_n8_n5# 0.07fF
C346 1bitaddie_3/ff_0/m1_106_n52# 1bitaddie_3/ff_0/m1_63_0# 0.05fF
C347 1bitaddie_0/sum 1bitaddie_0/xorg_1/m1_26_n95# 0.08fF
C348 vdd 1bitaddie_2/nandg_0/pmos_0/w_n8_n5# 0.08fF
C349 1bitaddie_2/inverter_1/out 1bitaddie_2/sum 0.20fF
C350 m1_560_235# ff_0/m1_106_n52# 0.05fF
C351 1bitaddie_2/ff_1/inverter_0/in vdd 0.12fF
C352 1bitaddie_2/xorg_0/pmos_1/w_n8_n5# 1bitaddie_2/xorg_0/m1_25_n11# 0.08fF
C353 1bitaddie_2/inverter_0/out 1bitaddie_2/Cin 0.02fF
C354 ff_1/inverter_0/in Cout 0.05fF
C355 1bitaddie_3/ff_1/pmos_1/w_n8_n5# 1bitaddie_3/ff_1/m1_19_n10# 0.08fF
C356 1bitaddie_2/inverter_0/w_n8_n5# 1bitaddie_2/inverter_0/in 0.07fF
C357 1bitaddie_2/xorg_0/inverter_1/w_n8_n5# 1bitaddie_2/xorg_0/inverter_1/out 0.03fF
C358 1bitaddie_2/ff_1/m1_106_n52# gnd 0.08fF
C359 1bitaddie_0/ff_2/m1_106_n52# gnd 0.08fF
C360 vdd s0 0.12fF
C361 1bitaddie_0/inverter_0/in 1bitaddie_0/Ai 0.13fF
C362 gnd 1bitaddie_1/xorg_0/inverter_1/out 0.08fF
C363 1bitaddie_4/xorg_1/pmos_2/w_n8_n5# vdd 0.08fF
C364 1bitaddie_0/ff_1/m1_63_0# vdd 0.12fF
C365 1bitaddie_0/xorg_0/inverter_0/w_n8_n5# 1bitaddie_0/xorg_0/inverter_0/out 0.03fF
C366 1bitaddie_2/ff_1/m1_58_n52# gnd 0.08fF
C367 1bitaddie_0/ff_2/m1_58_n52# gnd 0.08fF
C368 1bitaddie_4/manch_0/m1_24_n50# inverter_1/out 0.08fF
C369 1bitaddie_2/inverter_1/out 1bitaddie_4/clk 0.06fF
C370 1bitaddie_0/nandg_0/pmos_1/w_n8_n5# 1bitaddie_0/Ai 0.07fF
C371 1bitaddie_2/ff_0/m1_63_0# gnd 0.05fF
C372 1bitaddie_4/ff_0/m1_63_0# 1bitaddie_4/ff_0/pmos_3/w_n8_n5# 0.07fF
C373 1bitaddie_3/ff_1/inverter_0/in vdd 0.12fF
C374 1bitaddie_4/manch_0/clk 1bitaddie_4/Cin 0.07fF
C375 1bitaddie_2/inverter_0/out 1bitaddie_3/Cin 0.19fF
C376 1bitaddie_2/xorg_1/A 1bitaddie_2/xorg_1/m1_25_n11# 0.14fF
C377 1bitaddie_0/ff_1/m1_63_0# 1bitaddie_0/ff_1/m1_25_n37# 0.05fF
C378 1bitaddie_1/ff_1/inverter_0/in 1bitaddie_1/ff_1/m1_63_0# 0.05fF
C379 1bitaddie_1/ff_0/m1_58_n52# 1bitaddie_1/ff_0/m1_63_0# 0.08fF
C380 1bitaddie_4/ff_2/m1_63_0# gnd 0.05fF
C381 1bitaddie_3/ff_1/m1_106_n52# gnd 0.08fF
C382 1bitaddie_1/Bi 1bitaddie_1/inverter_0/in 0.11fF
C383 1bitaddie_3/inverter_0/out 1bitaddie_3/manch_0/clk 0.03fF
C384 1bitaddie_3/inverter_2/w_n8_n5# 1bitaddie_3/manch_0/clk 0.03fF
C385 1bitaddie_1/Ai 1bitaddie_1/nandg_0/m1_26_n48# 0.12fF
C386 1bitaddie_0/manch_0/clk vdd 0.12fF
C387 1bitaddie_4/inverter_2/w_n8_n5# 1bitaddie_4/clk 0.07fF
C388 1bitaddie_0/Ai 1bitaddie_0/xorg_0/m1_26_n95# 0.05fF
C389 m1_641_206# ff_0/pmos_1/w_n8_n5# 0.07fF
C390 1bitaddie_0/xorg_0/inverter_1/w_n8_n5# 1bitaddie_0/Bi 0.07fF
C391 1bitaddie_3/ff_1/m1_58_n52# gnd 0.08fF
C392 1bitaddie_3/inverter_1/out 1bitaddie_4/clk 0.06fF
C393 1bitaddie_1/ff_1/pmos_2/w_n8_n5# 1bitaddie_1/ff_1/m1_63_0# 0.03fF
C394 1bitaddie_2/ff_1/pmos_1/w_n8_n5# 1bitaddie_2/ff_1/m1_25_n37# 0.03fF
C395 1bitaddie_4/Bi 1bitaddie_4/clk 0.06fF
C396 1bitaddie_3/ff_0/m1_63_0# gnd 0.05fF
C397 1bitaddie_3/inverter_1/out 1bitaddie_3/sum 0.20fF
C398 1bitaddie_3/xorg_0/pmos_1/w_n8_n5# 1bitaddie_3/xorg_0/m1_25_n11# 0.08fF
C399 1bitaddie_0/ff_2/pmos_1/w_n8_n5# 1bitaddie_0/ff_2/m1_25_n37# 0.03fF
C400 1bitaddie_3/inverter_0/out 1bitaddie_3/Cin 0.02fF
C401 1bitaddie_4/inverter_1/out vdd 0.18fF
C402 1bitaddie_3/inverter_0/in 1bitaddie_3/nandg_0/m1_26_n48# 0.08fF
C403 1bitaddie_3/xorg_0/inverter_1/w_n8_n5# 1bitaddie_3/xorg_0/inverter_1/out 0.03fF
C404 vdd inverter_0/out 0.27fF
C405 1bitaddie_2/nandg_0/m1_26_n48# 1bitaddie_2/Ai 0.12fF
C406 1bitaddie_1/ff_0/inverter_0/in 1bitaddie_1/ff_0/m1_63_0# 0.05fF
C407 ff_0/m1_58_n52# ff_0/m1_63_0# 0.08fF
C408 1bitaddie_4/ff_0/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.07fF
C409 1bitaddie_1/ff_0/m1_63_0# 1bitaddie_1/ff_0/pmos_3/w_n8_n5# 0.07fF
C410 1bitaddie_1/xorg_0/inverter_1/out 1bitaddie_1/xorg_0/pmos_3/w_n8_n5# 0.07fF
C411 1bitaddie_1/xorg_0/pmos_0/w_n8_n5# 1bitaddie_1/xorg_0/m1_25_n11# 0.03fF
C412 1bitaddie_2/xorg_1/inverter_0/w_n8_n5# 1bitaddie_2/xorg_1/A 0.07fF
C413 1bitaddie_4/clk A1 0.17fF
C414 1bitaddie_0/ff_2/m1_63_0# 1bitaddie_0/ff_2/pmos_2/w_n8_n5# 0.03fF
C415 vdd 1bitaddie_1/ff_0/inverter_0/in 0.12fF
C416 1bitaddie_2/ff_2/m1_106_n52# gnd 0.08fF
C417 s2 vdd 0.12fF
C418 vdd 1bitaddie_1/ff_0/pmos_3/w_n8_n5# 0.06fF
C419 ff_1/pmos_0/w_n8_n5# ff_1/m1_19_n10# 0.03fF
C420 1bitaddie_3/xorg_1/A 1bitaddie_3/xorg_1/m1_25_n11# 0.14fF
C421 1bitaddie_4/Bi A4 0.03fF
C422 1bitaddie_4/inverter_1/w_n8_n5# vdd 0.08fF
C423 1bitaddie_4/clk 1bitaddie_1/ff_0/m1_25_n37# 0.31fF
C424 1bitaddie_4/ff_2/inverter_0/w_n8_n5# vdd 0.08fF
C425 vdd 1bitaddie_1/xorg_1/A 0.09fF
C426 inverter_1/out 1bitaddie_4/xorg_1/A 0.05fF
C427 1bitaddie_2/ff_1/m1_63_0# vdd 0.12fF
C428 1bitaddie_1/xorg_1/inverter_0/w_n8_n5# 1bitaddie_1/xorg_1/A 0.07fF
C429 1bitaddie_2/ff_2/m1_58_n52# gnd 0.08fF
C430 1bitaddie_2/xorg_1/pmos_3/w_n8_n5# 1bitaddie_2/xorg_1/m1_102_n17# 0.08fF
C431 1bitaddie_2/ff_2/pmos_1/w_n8_n5# 1bitaddie_2/ff_2/m1_19_n10# 0.08fF
C432 1bitaddie_2/Ai 1bitaddie_2/inverter_0/in 0.13fF
C433 1bitaddie_4/clk 1bitaddie_0/xorg_1/A 0.06fF
C434 1bitaddie_0/Bi 1bitaddie_0/ff_0/inverter_0/in 0.05fF
C435 1bitaddie_0/manch_0/pmos_0/w_n8_n5# 1bitaddie_1/Cin 0.03fF
C436 1bitaddie_3/ff_1/pmos_1/w_n8_n5# 1bitaddie_3/ff_1/m1_25_n37# 0.03fF
C437 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/sum 0.22fF
C438 gnd 1bitaddie_1/ff_0/m1_106_n52# 0.08fF
C439 1bitaddie_2/Bi 1bitaddie_2/ff_0/inverter_0/w_n8_n5# 0.03fF
C440 1bitaddie_1/ff_1/m1_25_n37# 1bitaddie_1/ff_1/m1_58_n52# 0.08fF
C441 1bitaddie_3/ff_2/m1_106_n52# gnd 0.08fF
C442 s3 vdd 0.12fF
C443 1bitaddie_3/inverter_1/w_n8_n5# vdd 0.08fF
C444 1bitaddie_0/inverter_0/out 1bitaddie_0/manch_0/m1_24_n50# 0.05fF
C445 1bitaddie_2/manch_0/clk vdd 0.12fF
C446 1bitaddie_0/xorg_0/pmos_2/w_n8_n5# 1bitaddie_0/xorg_0/m1_102_n17# 0.03fF
C447 1bitaddie_0/xorg_0/m1_26_n95# 1bitaddie_0/xorg_1/A 0.08fF
C448 1bitaddie_4/xorg_0/inverter_0/out 1bitaddie_4/clk 1.49fF
C449 1bitaddie_3/ff_1/m1_63_0# vdd 0.12fF
C450 1bitaddie_3/ff_2/m1_58_n52# gnd 0.08fF
C451 ff_1/m1_19_n10# vdd 0.12fF
C452 ff_1/m1_63_0# ff_1/m1_25_n37# 0.05fF
C453 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/xorg_1/pmos_3/w_n8_n5# 0.07fF
C454 1bitaddie_3/xorg_1/inverter_0/w_n8_n5# 1bitaddie_3/xorg_1/A 0.07fF
C455 1bitaddie_2/Cin vdd 0.12fF
C456 1bitaddie_4/clk 1bitaddie_1/ff_1/pmos_1/w_n8_n5# 0.31fF
C457 1bitaddie_0/xorg_1/pmos_0/w_n8_n5# 1bitaddie_0/xorg_1/m1_25_n11# 0.03fF
C458 1bitaddie_0/ff_2/inverter_0/in 1bitaddie_0/ff_2/m1_106_n52# 0.08fF
C459 1bitaddie_2/inverter_1/out 1bitaddie_2/xorg_1/pmos_1/w_n8_n5# 0.07fF
C460 1bitaddie_4/Ai vdd 0.21fF
C461 1bitaddie_2/sum 1bitaddie_2/xorg_1/m1_26_n95# 0.08fF
C462 1bitaddie_0/xorg_0/m1_102_n17# vdd 0.12fF
C463 1bitaddie_4/ff_1/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.07fF
C464 1bitaddie_3/manch_0/clk vdd 0.12fF
C465 1bitaddie_0/xorg_0/pmos_0/w_n8_n5# vdd 0.08fF
C466 1bitaddie_1/ff_1/pmos_0/w_n8_n5# 1bitaddie_1/ff_1/m1_19_n10# 0.03fF
C467 1bitaddie_3/xorg_1/pmos_3/w_n8_n5# 1bitaddie_3/xorg_1/m1_102_n17# 0.08fF
C468 1bitaddie_3/inverter_0/in 1bitaddie_3/Ai 0.13fF
C469 1bitaddie_4/xorg_0/inverter_1/out vdd 0.12fF
C470 1bitaddie_3/ff_2/pmos_1/w_n8_n5# 1bitaddie_3/ff_2/m1_19_n10# 0.08fF
C471 m1_560_235# ff_0/inverter_0/in 0.05fF
C472 vdd 1bitaddie_1/ff_1/m1_19_n10# 0.12fF
C473 vdd 1bitaddie_1/xorg_0/pmos_2/w_n8_n5# 0.08fF
C474 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/sum 0.22fF
C475 1bitaddie_3/Cin vdd 0.12fF
C476 1bitaddie_0/ff_2/inverter_0/in gnd 0.05fF
C477 ff_0/pmos_2/w_n8_n5# ff_0/m1_63_0# 0.03fF
C478 1bitaddie_3/Bi 1bitaddie_3/ff_0/inverter_0/w_n8_n5# 0.03fF
C479 1bitaddie_2/inverter_0/w_n8_n5# 1bitaddie_2/inverter_0/out 0.03fF
C480 1bitaddie_4/sum 1bitaddie_4/xorg_1/pmos_3/w_n8_n5# 0.03fF
C481 1bitaddie_4/xorg_1/inverter_1/out vdd 0.12fF
C482 1bitaddie_2/xorg_0/inverter_0/w_n8_n5# 1bitaddie_2/xorg_0/inverter_0/out 0.03fF
C483 1bitaddie_4/Ai 1bitaddie_4/ff_1/inverter_0/in 0.05fF
C484 1bitaddie_1/inverter_1/out 1bitaddie_1/xorg_1/A 0.06fF
C485 1bitaddie_1/ff_2/pmos_3/w_n8_n5# vdd 0.06fF
C486 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_4/clk 0.27fF
C487 1bitaddie_1/ff_0/inverter_0/w_n8_n5# 1bitaddie_1/ff_0/inverter_0/in 0.07fF
C488 1bitaddie_1/Bi 1bitaddie_1/xorg_0/inverter_1/out 0.05fF
C489 1bitaddie_2/xorg_1/A 1bitaddie_4/clk 0.06fF
C490 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_2/ff_1/m1_25_n37# 0.05fF
C491 1bitaddie_1/xorg_0/inverter_0/out 1bitaddie_4/clk 1.49fF
C492 ff_0/pmos_2/w_n8_n5# m1_608_244# 0.07fF
C493 1bitaddie_0/inverter_0/out 1bitaddie_0/xorg_1/A 0.06fF
C494 1bitaddie_0/ff_2/m1_63_0# 1bitaddie_0/ff_2/m1_106_n52# 0.05fF
C495 1bitaddie_2/Ai 1bitaddie_2/xorg_0/m1_26_n95# 0.05fF
C496 1bitaddie_0/xorg_1/pmos_2/w_n8_n5# vdd 0.08fF
C497 ff_0/pmos_1/w_n8_n5# ff_0/m1_25_n37# 0.03fF
C498 1bitaddie_4/ff_0/m1_106_n52# 1bitaddie_4/clk 0.05fF
C499 1bitaddie_2/xorg_0/inverter_1/w_n8_n5# 1bitaddie_2/Bi 0.07fF
C500 1bitaddie_3/inverter_1/out 1bitaddie_3/xorg_1/pmos_1/w_n8_n5# 0.07fF
C501 1bitaddie_4/xorg_1/inverter_0/out 1bitaddie_4/xorg_1/A 0.25fF
C502 1bitaddie_3/sum 1bitaddie_3/xorg_1/m1_26_n95# 0.08fF
C503 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_1/ff_2/m1_58_n52# 0.08fF
C504 gnd 1bitaddie_1/Bi 0.18fF
C505 1bitaddie_0/ff_2/m1_63_0# 1bitaddie_0/ff_2/m1_58_n52# 0.08fF
C506 1bitaddie_1/Ai vdd 0.21fF
C507 1bitaddie_4/ff_2/inverter_0/w_n8_n5# s4 0.03fF
C508 1bitaddie_2/ff_2/pmos_1/w_n8_n5# 1bitaddie_2/ff_2/m1_25_n37# 0.03fF
C509 1bitaddie_1/xorg_0/inverter_1/w_n8_n5# 1bitaddie_1/xorg_0/inverter_1/out 0.03fF
C510 1bitaddie_3/xorg_1/A 1bitaddie_4/clk 0.06fF
C511 1bitaddie_0/inverter_0/in 1bitaddie_0/Bi 0.11fF
C512 1bitaddie_4/clk 1bitaddie_1/ff_2/pmos_1/w_n8_n5# 0.07fF
C513 1bitaddie_0/ff_2/m1_63_0# gnd 0.05fF
C514 1bitaddie_4/clk B1 0.17fF
C515 1bitaddie_4/xorg_1/A vdd 0.09fF
C516 1bitaddie_4/inverter_0/in 1bitaddie_4/Ai 0.13fF
C517 1bitaddie_2/xorg_0/m1_102_n17# vdd 0.12fF
C518 1bitaddie_4/ff_2/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.28fF
C519 1bitaddie_2/xorg_0/pmos_0/w_n8_n5# vdd 0.08fF
C520 1bitaddie_4/clk 1bitaddie_0/inverter_2/w_n8_n5# 0.07fF
C521 1bitaddie_0/inverter_1/w_n8_n5# inverter_0/out 0.07fF
C522 1bitaddie_4/inverter_1/out 1bitaddie_4/Cin 0.05fF
C523 1bitaddie_3/xorg_0/inverter_0/w_n8_n5# 1bitaddie_3/xorg_0/inverter_0/out 0.03fF
C524 1bitaddie_1/ff_2/pmos_3/w_n8_n5# 1bitaddie_1/ff_2/inverter_0/in 0.03fF
C525 1bitaddie_2/ff_2/m1_63_0# 1bitaddie_2/ff_2/pmos_2/w_n8_n5# 0.03fF
C526 1bitaddie_4/clk 1bitaddie_1/ff_1/m1_63_0# 0.35fF
C527 B4 gnd 0.05fF
C528 1bitaddie_4/ff_0/inverter_0/in gnd 0.05fF
C529 1bitaddie_4/xorg_0/inverter_1/out 1bitaddie_4/xorg_0/m1_102_n91# 0.05fF
C530 1bitaddie_4/clk 1bitaddie_0/Bi 0.06fF
C531 1bitaddie_0/ff_1/m1_63_0# 1bitaddie_0/ff_1/inverter_0/in 0.05fF
C532 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_3/ff_1/m1_25_n37# 0.05fF
C533 vdd 1bitaddie_1/ff_2/m1_19_n10# 0.12fF
C534 1bitaddie_4/inverter_0/w_n8_n5# vdd 0.08fF
C535 1bitaddie_0/inverter_1/out vdd 0.18fF
C536 1bitaddie_2/ff_2/inverter_0/in gnd 0.05fF
C537 1bitaddie_1/nandg_0/pmos_1/w_n8_n5# 1bitaddie_1/inverter_0/in 0.03fF
C538 ff_0/m1_63_0# vdd 0.12fF
C539 1bitaddie_0/Bi 1bitaddie_0/xorg_0/m1_26_n95# 0.05fF
C540 1bitaddie_3/xorg_0/m1_102_n17# vdd 0.12fF
C541 1bitaddie_4/clk 1bitaddie_0/ff_0/pmos_2/w_n8_n5# 0.07fF
C542 1bitaddie_0/ff_0/inverter_0/in 1bitaddie_0/ff_0/m1_106_n52# 0.08fF
C543 1bitaddie_3/xorg_0/pmos_0/w_n8_n5# vdd 0.08fF
C544 1bitaddie_3/Ai 1bitaddie_3/xorg_0/m1_26_n95# 0.05fF
C545 1bitaddie_3/xorg_0/inverter_1/w_n8_n5# 1bitaddie_3/Bi 0.07fF
C546 1bitaddie_4/clk 1bitaddie_1/ff_0/pmos_1/w_n8_n5# 0.30fF
C547 1bitaddie_4/clk 1bitaddie_1/inverter_2/w_n8_n5# 0.07fF
C548 ff_0/pmos_0/w_n8_n5# C0 0.07fF
C549 1bitaddie_4/ff_1/m1_106_n52# 1bitaddie_4/clk 0.05fF
C550 1bitaddie_4/inverter_1/w_n8_n5# 1bitaddie_4/Cin 0.07fF
C551 1bitaddie_2/Bi 1bitaddie_2/ff_0/inverter_0/in 0.05fF
C552 vdd 1bitaddie_2/nandg_0/pmos_1/w_n8_n5# 0.08fF
C553 1bitaddie_4/sum gnd 0.35fF
C554 1bitaddie_4/nandg_0/pmos_0/w_n8_n5# 1bitaddie_4/Bi 0.07fF
C555 1bitaddie_0/sum 1bitaddie_0/xorg_1/m1_102_n17# 0.12fF
C556 1bitaddie_3/ff_2/pmos_1/w_n8_n5# 1bitaddie_3/ff_2/m1_25_n37# 0.03fF
C557 1bitaddie_2/nandg_0/m1_26_n48# 1bitaddie_2/Bi 0.05fF
C558 1bitaddie_2/inverter_0/out 1bitaddie_2/manch_0/m1_24_n50# 0.05fF
C559 1bitaddie_2/xorg_0/pmos_2/w_n8_n5# 1bitaddie_2/xorg_0/m1_102_n17# 0.03fF
C560 1bitaddie_2/xorg_0/m1_26_n95# 1bitaddie_2/xorg_1/A 0.08fF
C561 1bitaddie_4/ff_1/m1_58_n52# 1bitaddie_4/clk 0.12fF
C562 1bitaddie_3/ff_2/inverter_0/in gnd 0.05fF
C563 1bitaddie_2/xorg_1/pmos_2/w_n8_n5# vdd 0.08fF
C564 1bitaddie_1/inverter_0/out 1bitaddie_1/Cin 0.02fF
C565 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/xorg_1/m1_102_n91# 0.05fF
C566 1bitaddie_0/ff_2/inverter_0/w_n8_n5# vdd 0.08fF
C567 1bitaddie_4/ff_0/m1_63_0# 1bitaddie_4/clk 0.35fF
C568 ff_1/inverter_0/w_n8_n5# ff_1/inverter_0/in 0.07fF
C569 vdd 1bitaddie_1/ff_0/m1_19_n10# 0.12fF
C570 1bitaddie_4/ff_0/inverter_0/w_n8_n5# 1bitaddie_4/ff_0/inverter_0/in 0.07fF
C571 1bitaddie_3/ff_2/m1_63_0# 1bitaddie_3/ff_2/pmos_2/w_n8_n5# 0.03fF
C572 1bitaddie_1/xorg_0/m1_26_n95# 1bitaddie_1/xorg_1/A 0.08fF
C573 1bitaddie_2/xorg_1/pmos_0/w_n8_n5# 1bitaddie_2/xorg_1/m1_25_n11# 0.03fF
C574 1bitaddie_2/ff_2/m1_63_0# gnd 0.05fF
C575 1bitaddie_2/ff_2/inverter_0/in 1bitaddie_2/ff_2/m1_106_n52# 0.08fF
C576 1bitaddie_1/ff_2/pmos_3/w_n8_n5# 1bitaddie_1/ff_2/m1_63_0# 0.07fF
C577 1bitaddie_4/manch_0/m1_24_n50# 1bitaddie_4/manch_0/clk 0.05fF
C578 1bitaddie_4/xorg_0/m1_102_n91# 1bitaddie_4/xorg_1/A 0.08fF
C579 1bitaddie_0/Ai 1bitaddie_0/xorg_0/pmos_2/w_n8_n5# 0.07fF
C580 1bitaddie_3/xorg_1/pmos_2/w_n8_n5# vdd 0.08fF
C581 1bitaddie_2/Bi 1bitaddie_2/inverter_0/in 0.11fF
C582 1bitaddie_4/clk 1bitaddie_0/xorg_0/inverter_0/out 1.49fF
C583 1bitaddie_2/inverter_0/w_n8_n5# vdd 0.08fF
C584 1bitaddie_1/ff_2/pmos_0/w_n8_n5# 1bitaddie_1/ff_2/m1_19_n10# 0.03fF
C585 ff_0/m1_106_n52# gnd 0.08fF
C586 1bitaddie_2/Bi 1bitaddie_4/clk 0.06fF
C587 1bitaddie_4/clk 1bitaddie_1/Cin 0.11fF
C588 1bitaddie_3/Bi 1bitaddie_3/ff_0/inverter_0/in 0.05fF
C589 1bitaddie_3/manch_0/clk 1bitaddie_4/Cin 0.16fF
C590 1bitaddie_4/manch_0/m1_24_n50# 1bitaddie_4/Cin 0.07fF
C591 1bitaddie_2/inverter_1/out vdd 0.18fF
C592 1bitaddie_4/inverter_0/in 1bitaddie_4/inverter_0/w_n8_n5# 0.07fF
C593 1bitaddie_3/ff_2/m1_63_0# gnd 0.05fF
C594 1bitaddie_4/ff_0/m1_63_0# 1bitaddie_4/ff_0/m1_25_n37# 0.05fF
C595 1bitaddie_3/inverter_0/out 1bitaddie_3/manch_0/m1_24_n50# 0.05fF
C596 1bitaddie_3/xorg_0/pmos_2/w_n8_n5# 1bitaddie_3/xorg_0/m1_102_n17# 0.03fF
C597 1bitaddie_0/xorg_1/m1_102_n91# 1bitaddie_0/xorg_1/inverter_0/out 0.05fF
C598 1bitaddie_0/Ai vdd 0.21fF
C599 1bitaddie_3/xorg_0/m1_26_n95# 1bitaddie_3/xorg_1/A 0.08fF
C600 1bitaddie_2/ff_0/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.07fF
C601 1bitaddie_1/xorg_1/m1_26_n95# 1bitaddie_1/sum 0.08fF
C602 1bitaddie_4/clk 1bitaddie_0/ff_1/pmos_2/w_n8_n5# 0.07fF
C603 1bitaddie_0/ff_0/inverter_0/in 1bitaddie_0/ff_0/m1_63_0# 0.05fF
C604 1bitaddie_4/ff_2/m1_106_n52# 1bitaddie_4/clk 0.05fF
C605 1bitaddie_3/Cin 1bitaddie_4/Cin 0.14fF
C606 1bitaddie_1/xorg_1/A 1bitaddie_1/xorg_1/m1_102_n17# 0.20fF
C607 1bitaddie_1/inverter_0/out 1bitaddie_1/inverter_0/in 0.05fF
C608 1bitaddie_0/xorg_0/inverter_1/out vdd 0.12fF
C609 1bitaddie_4/inverter_2/w_n8_n5# vdd 0.08fF
C610 1bitaddie_3/Bi 1bitaddie_4/clk 0.06fF
C611 1bitaddie_2/inverter_0/out 1bitaddie_2/xorg_1/A 0.06fF
C612 1bitaddie_2/ff_2/m1_63_0# 1bitaddie_2/ff_2/m1_106_n52# 0.05fF
C613 1bitaddie_4/clk 1bitaddie_1/sum 0.08fF
C614 inverter_0/in vdd 0.12fF
C615 1bitaddie_3/inverter_1/out vdd 0.18fF
C616 1bitaddie_3/xorg_1/pmos_0/w_n8_n5# 1bitaddie_3/xorg_1/m1_25_n11# 0.03fF
C617 1bitaddie_1/manch_0/clk 1bitaddie_2/Cin 0.16fF
C618 1bitaddie_4/ff_2/m1_58_n52# 1bitaddie_4/clk 0.11fF
C619 1bitaddie_4/Bi vdd 0.24fF
C620 1bitaddie_3/ff_2/inverter_0/in 1bitaddie_3/ff_2/m1_106_n52# 0.08fF
C621 gnd 1bitaddie_1/ff_1/inverter_0/in 0.05fF
C622 1bitaddie_0/ff_2/inverter_0/in 1bitaddie_0/ff_2/m1_63_0# 0.05fF
C623 1bitaddie_2/ff_2/inverter_0/w_n8_n5# vdd 0.08fF
C624 ff_0/m1_19_n10# ff_0/m1_25_n37# 0.12fF
C625 vdd 1bitaddie_1/xorg_1/inverter_0/out 0.12fF
C626 1bitaddie_0/xorg_1/inverter_1/out vdd 0.12fF
C627 1bitaddie_2/ff_2/m1_63_0# 1bitaddie_2/ff_2/m1_58_n52# 0.08fF
C628 1bitaddie_3/ff_0/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.07fF
C629 1bitaddie_1/ff_1/m1_63_0# 1bitaddie_1/ff_1/m1_106_n52# 0.05fF
C630 1bitaddie_1/xorg_1/inverter_0/w_n8_n5# 1bitaddie_1/xorg_1/inverter_0/out 0.03fF
C631 1bitaddie_3/inverter_0/in 1bitaddie_3/Bi 0.11fF
C632 1bitaddie_4/sum 1bitaddie_4/xorg_1/m1_25_n11# 0.12fF
C633 1bitaddie_1/ff_1/pmos_0/w_n8_n5# A1 0.07fF
C634 1bitaddie_4/ff_0/pmos_2/w_n8_n5# vdd 0.08fF
C635 1bitaddie_1/ff_1/m1_63_0# 1bitaddie_1/ff_1/m1_58_n52# 0.08fF
C636 1bitaddie_1/ff_0/m1_63_0# 1bitaddie_1/ff_0/m1_25_n37# 0.05fF
C637 1bitaddie_4/xorg_0/m1_26_n95# gnd 0.08fF
C638 inverter_1/in ff_1/m1_19_n10# 0.11fF
C639 1bitaddie_4/clk 1bitaddie_2/inverter_2/w_n8_n5# 0.07fF
C640 1bitaddie_3/ff_2/inverter_0/w_n8_n5# vdd 0.08fF
C641 1bitaddie_4/clk 1bitaddie_0/ff_0/m1_106_n52# 0.05fF
C642 1bitaddie_2/xorg_0/inverter_0/out 1bitaddie_4/clk 1.49fF
C643 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_2/ff_1/inverter_0/in 0.05fF
C644 1bitaddie_4/xorg_1/A 1bitaddie_4/Cin 0.10fF
C645 1bitaddie_0/ff_0/m1_63_0# 1bitaddie_0/ff_0/pmos_3/w_n8_n5# 0.07fF
C646 1bitaddie_0/manch_0/clk inverter_0/out 0.07fF
C647 1bitaddie_0/inverter_0/out 1bitaddie_1/Cin 0.19fF
C648 1bitaddie_4/ff_1/m1_58_n52# 1bitaddie_4/ff_1/m1_25_n37# 0.08fF
C649 ff_1/inverter_0/in gnd 0.05fF
C650 ff_0/m1_63_0# ff_0/pmos_3/w_n8_n5# 0.07fF
C651 1bitaddie_4/ff_2/inverter_0/in 1bitaddie_4/ff_2/pmos_3/w_n8_n5# 0.03fF
C652 1bitaddie_4/Ai 1bitaddie_4/xorg_0/m1_102_n17# 0.20fF
C653 1bitaddie_3/inverter_0/out 1bitaddie_3/xorg_1/A 0.06fF
C654 1bitaddie_3/ff_2/m1_63_0# 1bitaddie_3/ff_2/m1_106_n52# 0.05fF
C655 1bitaddie_2/Bi 1bitaddie_2/xorg_0/m1_26_n95# 0.05fF
C656 1bitaddie_1/Ai 1bitaddie_1/xorg_0/m1_26_n95# 0.05fF
C657 1bitaddie_2/ff_0/inverter_0/in 1bitaddie_2/ff_0/m1_106_n52# 0.08fF
C658 1bitaddie_1/xorg_0/inverter_1/w_n8_n5# 1bitaddie_1/Bi 0.07fF
C659 1bitaddie_0/xorg_1/A vdd 0.09fF
C660 1bitaddie_2/Ai vdd 0.21fF
C661 1bitaddie_0/inverter_1/w_n8_n5# 1bitaddie_0/inverter_1/out 0.03fF
C662 1bitaddie_4/sum 1bitaddie_4/ff_2/pmos_0/w_n8_n5# 0.07fF
C663 1bitaddie_2/ff_1/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.07fF
C664 1bitaddie_4/clk 1bitaddie_0/ff_2/pmos_2/w_n8_n5# 0.28fF
C665 1bitaddie_3/xorg_0/inverter_0/out 1bitaddie_4/clk 1.49fF
C666 1bitaddie_3/ff_2/m1_63_0# 1bitaddie_3/ff_2/m1_58_n52# 0.08fF
C667 B0 gnd 0.05fF
C668 1bitaddie_2/sum 1bitaddie_2/xorg_1/m1_102_n17# 0.12fF
C669 1bitaddie_2/xorg_0/inverter_1/out vdd 0.12fF
C670 1bitaddie_1/manch_0/m1_24_n50# 1bitaddie_1/manch_0/clk 0.05fF
C671 1bitaddie_0/ff_0/inverter_0/in gnd 0.05fF
C672 1bitaddie_4/xorg_0/inverter_0/out vdd 0.12fF
C673 1bitaddie_3/inverter_0/in 1bitaddie_3/nandg_0/pmos_0/w_n8_n5# 0.03fF
C674 vdd 1bitaddie_1/xorg_1/m1_25_n11# 0.12fF
C675 1bitaddie_4/inverter_0/in 1bitaddie_4/Bi 0.11fF
C676 1bitaddie_4/xorg_0/m1_25_n11# vdd 0.12fF
C677 1bitaddie_2/xorg_1/inverter_1/out vdd 0.12fF
C678 1bitaddie_3/Ai vdd 0.21fF
C679 1bitaddie_3/ff_1/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.07fF
C680 1bitaddie_4/inverter_1/w_n8_n5# 1bitaddie_4/inverter_1/out 0.03fF
C681 1bitaddie_4/clk 1bitaddie_0/ff_1/m1_106_n52# 0.05fF
C682 1bitaddie_4/ff_1/pmos_2/w_n8_n5# vdd 0.08fF
C683 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/xorg_1/m1_102_n91# 0.05fF
C684 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_3/ff_1/inverter_0/in 0.05fF
C685 1bitaddie_3/xorg_0/inverter_1/out vdd 0.12fF
C686 1bitaddie_0/sum gnd 0.35fF
C687 ff_1/m1_106_n52# gnd 0.08fF
C688 Cout vdd 0.12fF
C689 1bitaddie_4/inverter_0/out gnd 0.08fF
C690 1bitaddie_4/ff_2/m1_63_0# 1bitaddie_4/ff_2/pmos_3/w_n8_n5# 0.07fF
C691 1bitaddie_4/inverter_0/in 1bitaddie_4/nandg_0/m1_26_n48# 0.08fF
C692 1bitaddie_2/Ai 1bitaddie_2/xorg_0/pmos_2/w_n8_n5# 0.07fF
C693 1bitaddie_4/clk 1bitaddie_0/ff_1/m1_58_n52# 0.12fF
C694 1bitaddie_3/Bi 1bitaddie_3/xorg_0/m1_26_n95# 0.05fF
C695 1bitaddie_1/ff_0/inverter_0/in 1bitaddie_1/ff_0/pmos_3/w_n8_n5# 0.03fF
C696 1bitaddie_0/Bi A0 0.03fF
C697 m1_641_206# ff_0/m1_25_n37# 0.06fF
C698 1bitaddie_2/ff_0/m1_106_n52# 1bitaddie_4/clk 0.05fF
C699 ff_1/m1_58_n52# gnd 0.08fF
C700 1bitaddie_3/ff_0/inverter_0/in 1bitaddie_3/ff_0/m1_106_n52# 0.08fF
C701 1bitaddie_3/xorg_1/inverter_1/out vdd 0.12fF
C702 1bitaddie_4/clk 1bitaddie_0/ff_0/m1_63_0# 0.35fF
C703 1bitaddie_4/xorg_1/inverter_0/out 1bitaddie_4/xorg_1/pmos_0/w_n8_n5# 0.07fF
C704 1bitaddie_0/inverter_0/in 1bitaddie_0/nandg_0/pmos_0/w_n8_n5# 0.03fF
C705 ff_0/inverter_0/in gnd 0.05fF
C706 1bitaddie_1/xorg_1/pmos_3/w_n8_n5# 1bitaddie_1/xorg_1/m1_102_n17# 0.08fF
C707 1bitaddie_3/sum 1bitaddie_3/xorg_1/m1_102_n17# 0.12fF
C708 1bitaddie_4/xorg_0/m1_102_n17# 1bitaddie_4/xorg_1/A 0.12fF
C709 1bitaddie_4/xorg_1/m1_102_n17# vdd 0.12fF
C710 1bitaddie_2/xorg_1/m1_102_n91# 1bitaddie_2/xorg_1/inverter_0/out 0.05fF
C711 1bitaddie_1/xorg_0/inverter_0/out vdd 0.12fF
C712 1bitaddie_4/ff_0/m1_63_0# 1bitaddie_4/ff_0/m1_58_n52# 0.08fF
C713 1bitaddie_4/xorg_1/pmos_0/w_n8_n5# vdd 0.08fF
C714 1bitaddie_2/xorg_1/A vdd 0.09fF
C715 inverter_1/in ff_1/m1_25_n37# 0.05fF
C716 1bitaddie_2/ff_2/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.28fF
C717 1bitaddie_2/ff_0/inverter_0/in 1bitaddie_2/ff_0/m1_63_0# 0.05fF
C718 1bitaddie_1/nandg_0/pmos_0/w_n8_n5# vdd 0.08fF
C719 1bitaddie_3/ff_0/m1_106_n52# 1bitaddie_4/clk 0.05fF
C720 1bitaddie_4/inverter_2/w_n8_n5# 1bitaddie_4/manch_0/clk 0.03fF
C721 1bitaddie_4/xorg_0/pmos_3/w_n8_n5# 1bitaddie_4/xorg_0/m1_102_n17# 0.08fF
C722 B2 gnd 0.05fF
C723 1bitaddie_4/ff_0/inverter_0/in 1bitaddie_4/ff_0/pmos_3/w_n8_n5# 0.03fF
C724 1bitaddie_2/ff_0/inverter_0/in gnd 0.05fF
C725 1bitaddie_4/ff_2/inverter_0/in 1bitaddie_4/clk 0.05fF
C726 1bitaddie_4/xorg_0/inverter_0/out 1bitaddie_4/xorg_0/m1_102_n91# 0.05fF
C727 1bitaddie_2/ff_2/inverter_0/in 1bitaddie_2/ff_2/m1_63_0# 0.05fF
C728 1bitaddie_2/nandg_0/m1_26_n48# gnd 0.08fF
C729 1bitaddie_1/inverter_0/out gnd 0.08fF
C730 1bitaddie_1/inverter_0/in 1bitaddie_1/nandg_0/m1_26_n48# 0.08fF
C731 1bitaddie_3/xorg_1/A vdd 0.09fF
C732 1bitaddie_3/Ai 1bitaddie_3/xorg_0/pmos_2/w_n8_n5# 0.07fF
C733 1bitaddie_4/xorg_1/pmos_1/w_n8_n5# 1bitaddie_4/xorg_1/m1_25_n11# 0.08fF
C734 1bitaddie_3/ff_2/pmos_2/w_n8_n5# 1bitaddie_4/clk 0.28fF
C735 1bitaddie_2/ff_1/m1_106_n52# 1bitaddie_4/clk 0.05fF
C736 1bitaddie_4/clk 1bitaddie_0/ff_2/m1_106_n52# 0.05fF
C737 1bitaddie_4/ff_2/pmos_2/w_n8_n5# vdd 0.08fF
C738 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/inverter_1/out 0.05fF
C739 B3 gnd 0.05fF
C740 1bitaddie_2/sum gnd 0.35fF
C741 1bitaddie_2/Cin 1bitaddie_1/xorg_1/A 0.05fF
C742 1bitaddie_3/ff_0/inverter_0/in gnd 0.05fF
C743 1bitaddie_0/inverter_2/w_n8_n5# vdd 0.08fF
C744 1bitaddie_0/inverter_0/in gnd 0.05fF
C745 1bitaddie_4/xorg_1/A 1bitaddie_4/xorg_1/pmos_2/w_n8_n5# 0.07fF
C746 1bitaddie_4/xorg_1/inverter_1/w_n8_n5# vdd 0.08fF
C747 vdd 1bitaddie_1/ff_1/m1_63_0# 0.12fF
C748 1bitaddie_2/ff_1/m1_58_n52# 1bitaddie_4/clk 0.12fF
C749 vdd 1bitaddie_2/inverter_1/w_n8_n5# 0.08fF
C750 1bitaddie_1/xorg_1/m1_26_n95# gnd 0.08fF
C751 1bitaddie_4/clk 1bitaddie_0/ff_2/m1_58_n52# 0.11fF
C752 1bitaddie_0/Bi vdd 0.24fF
C753 1bitaddie_3/xorg_1/m1_102_n91# 1bitaddie_3/xorg_1/inverter_0/out 0.05fF
C754 m1_611_197# ff_0/m1_25_n37# 0.07fF
C755 1bitaddie_2/ff_0/m1_63_0# 1bitaddie_4/clk 0.35fF
C756 1bitaddie_0/sum 1bitaddie_0/xorg_1/pmos_3/w_n8_n5# 0.03fF
C757 1bitaddie_3/ff_0/inverter_0/in 1bitaddie_3/ff_0/m1_63_0# 0.05fF
C758 gnd 1bitaddie_2/inverter_0/in 0.05fF
C759 vdd 1bitaddie_1/ff_0/pmos_0/w_n8_n5# 0.08fF
C760 1bitaddie_0/Ai 1bitaddie_0/ff_1/inverter_0/in 0.05fF
C761 1bitaddie_2/ff_0/m1_63_0# 1bitaddie_2/ff_0/pmos_3/w_n8_n5# 0.07fF
C762 1bitaddie_4/ff_2/m1_63_0# 1bitaddie_4/clk 0.27fF
C763 1bitaddie_3/ff_1/m1_106_n52# 1bitaddie_4/clk 0.05fF
C764 1bitaddie_2/manch_0/clk 1bitaddie_2/Cin 0.07fF
C765 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/sum 0.22fF
C766 1bitaddie_4/clk gnd 2.60fF
C767 1bitaddie_0/ff_0/pmos_2/w_n8_n5# vdd 0.08fF
C768 1bitaddie_3/sum gnd 0.35fF
C769 1bitaddie_4/ff_2/m1_58_n52# 1bitaddie_4/ff_2/m1_25_n37# 0.08fF
C770 vdd 1bitaddie_1/inverter_2/w_n8_n5# 0.08fF
C771 gnd 1bitaddie_1/ff_2/m1_106_n52# 0.08fF
C772 vdd s1 0.12fF
C773 1bitaddie_0/xorg_0/m1_26_n95# gnd 0.08fF
C774 1bitaddie_4/inverter_1/out 1bitaddie_4/xorg_1/m1_26_n95# 0.05fF
C775 1bitaddie_3/ff_2/inverter_0/in 1bitaddie_3/ff_2/m1_63_0# 0.05fF
C776 1bitaddie_3/ff_1/m1_58_n52# 1bitaddie_4/clk 0.12fF
C777 1bitaddie_3/ff_0/m1_63_0# 1bitaddie_4/clk 0.35fF
C778 1bitaddie_3/inverter_0/in gnd 0.05fF
C779 1bitaddie_0/xorg_1/inverter_0/out 1bitaddie_0/xorg_1/A 0.25fF
C780 1bitaddie_4/inverter_1/out 1bitaddie_4/xorg_1/A 0.06fF
C781 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/ff_1/pmos_2/w_n8_n5# 0.03fF
C782 gnd 1bitaddie_1/ff_2/m1_58_n52# 0.08fF
C783 1bitaddie_3/inverter_1/w_n8_n5# 1bitaddie_3/Cin 0.07fF
C784 1bitaddie_0/ff_2/inverter_0/w_n8_n5# s0 0.03fF
C785 1bitaddie_4/ff_0/m1_63_0# vdd 0.12fF
C786 1bitaddie_2/manch_0/clk 1bitaddie_3/Cin 0.16fF
C787 A4 gnd 0.05fF
C788 1bitaddie_4/ff_1/inverter_0/in 1bitaddie_4/ff_1/m1_106_n52# 0.08fF
C789 1bitaddie_3/nandg_0/pmos_1/w_n8_n5# 1bitaddie_3/Ai 0.07fF
C790 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_1/ff_2/m1_63_0# 0.05fF
C791 1bitaddie_4/ff_0/m1_25_n37# gnd 0.08fF
C792 1bitaddie_2/Cin 1bitaddie_3/Cin 0.14fF
C793 1bitaddie_0/inverter_1/out inverter_0/out 0.05fF
C794 1bitaddie_2/ff_2/m1_106_n52# 1bitaddie_4/clk 0.05fF
C795 1bitaddie_0/xorg_0/inverter_1/out 1bitaddie_0/xorg_0/m1_102_n91# 0.05fF
C796 1bitaddie_4/Bi 1bitaddie_4/xorg_0/m1_102_n17# 0.05fF
C797 1bitaddie_3/ff_0/m1_63_0# 1bitaddie_3/ff_0/pmos_3/w_n8_n5# 0.07fF
C798 1bitaddie_0/xorg_0/inverter_0/out vdd 0.12fF
C799 1bitaddie_3/manch_0/clk 1bitaddie_3/Cin 0.07fF
C800 1bitaddie_3/manch_0/m1_24_n50# 1bitaddie_4/Cin 0.08fF
C801 1bitaddie_2/Bi A2 0.03fF
C802 1bitaddie_2/Bi vdd 0.24fF
C803 s1 1bitaddie_1/ff_2/inverter_0/in 0.05fF
C804 vdd 1bitaddie_1/Cin 0.12fF
C805 1bitaddie_2/ff_2/m1_58_n52# 1bitaddie_4/clk 0.11fF
C806 ff_0/inverter_0/in ff_0/inverter_0/w_n8_n5# 0.07fF
C807 1bitaddie_1/inverter_0/out 1bitaddie_1/inverter_0/w_n8_n5# 0.03fF
C808 1bitaddie_0/xorg_0/m1_25_n11# vdd 0.12fF
C809 1bitaddie_4/clk 1bitaddie_1/ff_0/m1_106_n52# 0.05fF
C810 1bitaddie_3/ff_2/m1_106_n52# 1bitaddie_4/clk 0.05fF
C811 1bitaddie_2/ff_0/pmos_2/w_n8_n5# vdd 0.08fF
C812 1bitaddie_0/ff_1/pmos_2/w_n8_n5# vdd 0.08fF
C813 vdd 1bitaddie_1/xorg_0/m1_102_n17# 0.12fF
C814 vdd 1bitaddie_1/xorg_0/pmos_0/w_n8_n5# 0.08fF
C815 1bitaddie_0/inverter_0/out gnd 0.08fF
C816 1bitaddie_4/ff_1/pmos_0/w_n8_n5# 1bitaddie_4/ff_1/m1_19_n10# 0.03fF
C817 1bitaddie_2/xorg_0/m1_26_n95# gnd 0.08fF
C818 1bitaddie_3/Bi vdd 0.24fF
C819 1bitaddie_1/manch_0/m1_24_n50# 1bitaddie_2/Cin 0.08fF
C820 1bitaddie_4/sum 1bitaddie_4/xorg_1/pmos_1/w_n8_n5# 0.03fF
C821 1bitaddie_3/ff_2/m1_58_n52# 1bitaddie_4/clk 0.11fF
C822 1bitaddie_0/inverter_0/w_n8_n5# 1bitaddie_0/inverter_0/in 0.07fF
C823 A4 1bitaddie_4/ff_1/pmos_0/w_n8_n5# 0.07fF
C824 1bitaddie_0/ff_0/inverter_0/w_n8_n5# 1bitaddie_0/ff_0/inverter_0/in 0.07fF
C825 1bitaddie_3/ff_0/pmos_2/w_n8_n5# vdd 0.08fF
C826 1bitaddie_1/Ai 1bitaddie_1/xorg_0/pmos_2/w_n8_n5# 0.07fF
C827 ff_1/m1_19_n10# ff_1/m1_25_n37# 0.12fF
C828 ff_0/m1_58_n52# gnd 0.08fF
C829 1bitaddie_0/xorg_1/m1_102_n17# vdd 0.12fF
C830 1bitaddie_3/xorg_0/m1_26_n95# gnd 0.08fF
C831 1bitaddie_3/Bi A3 0.03fF
C832 1bitaddie_0/xorg_1/pmos_0/w_n8_n5# vdd 0.08fF
C833 1bitaddie_0/manch_0/m1_24_n50# 1bitaddie_0/manch_0/clk 0.05fF
C834 1bitaddie_0/xorg_0/m1_102_n91# 1bitaddie_0/xorg_1/A 0.08fF
C835 1bitaddie_4/xorg_0/inverter_1/out 1bitaddie_4/xorg_1/A 0.22fF
C836 1bitaddie_4/ff_1/m1_25_n37# gnd 0.08fF
C837 vdd 1bitaddie_2/inverter_2/w_n8_n5# 0.08fF
C838 gnd 1bitaddie_1/ff_1/m1_106_n52# 0.08fF
C839 1bitaddie_4/xorg_0/inverter_0/out 1bitaddie_4/xorg_0/pmos_0/w_n8_n5# 0.07fF
C840 vdd 1bitaddie_1/inverter_0/in 0.25fF
C841 gnd 1bitaddie_1/nandg_0/m1_26_n48# 0.08fF
C842 1bitaddie_3/xorg_1/A 1bitaddie_4/Cin 0.05fF
C843 1bitaddie_2/xorg_0/inverter_0/out vdd 0.12fF
C844 1bitaddie_4/clk 1bitaddie_0/ff_2/inverter_0/in 0.05fF
C845 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/ff_1/m1_106_n52# 0.05fF
C846 1bitaddie_4/xorg_0/inverter_1/out 1bitaddie_4/xorg_0/pmos_3/w_n8_n5# 0.07fF
C847 1bitaddie_4/xorg_0/pmos_0/w_n8_n5# 1bitaddie_4/xorg_0/m1_25_n11# 0.03fF
C848 1bitaddie_0/manch_0/m1_24_n50# inverter_0/out 0.07fF
C849 B4 1bitaddie_4/ff_0/m1_19_n10# 0.11fF
C850 gnd 1bitaddie_1/ff_1/m1_58_n52# 0.08fF
C851 1bitaddie_2/xorg_0/m1_25_n11# vdd 0.12fF
C852 1bitaddie_2/sum 1bitaddie_2/xorg_1/pmos_3/w_n8_n5# 0.03fF
C853 ff_1/nmos_2/a_0_n10# ff_1/m1_25_n37# 0.03fF
C854 1bitaddie_0/ff_0/m1_63_0# 1bitaddie_0/ff_0/m1_25_n37# 0.05fF
C855 1bitaddie_1/Cin 1bitaddie_1/inverter_1/out 0.05fF
C856 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/ff_1/m1_58_n52# 0.08fF
C857 1bitaddie_2/Ai 1bitaddie_2/ff_1/inverter_0/in 0.05fF
C858 ff_0/m1_63_0# ff_0/m1_25_n37# 0.05fF
C859 1bitaddie_3/nandg_0/pmos_0/w_n8_n5# vdd 0.08fF
C860 inverter_0/in inverter_0/out 0.05fF
C861 1bitaddie_2/ff_1/pmos_2/w_n8_n5# vdd 0.08fF
C862 vdd 1bitaddie_0/ff_2/pmos_2/w_n8_n5# 0.08fF
C863 1bitaddie_3/xorg_0/inverter_0/out vdd 0.12fF
C864 1bitaddie_2/inverter_0/out gnd 0.08fF
C865 1bitaddie_1/ff_2/pmos_0/w_n8_n5# 1bitaddie_1/sum 0.07fF
C866 1bitaddie_0/xorg_1/inverter_1/w_n8_n5# vdd 0.08fF
C867 1bitaddie_3/xorg_0/m1_25_n11# vdd 0.12fF
C868 1bitaddie_4/clk 1bitaddie_1/Bi 0.06fF
C869 inverter_1/out gnd 0.12fF
C870 1bitaddie_4/xorg_1/m1_26_n95# 1bitaddie_4/xorg_1/A 0.05fF
C871 1bitaddie_2/xorg_1/inverter_0/out 1bitaddie_2/xorg_1/A 0.25fF
C872 1bitaddie_1/ff_1/m1_19_n10# 1bitaddie_1/ff_1/m1_25_n37# 0.12fF
C873 ff_1/inverter_0/w_n8_n5# vdd 0.08fF
C874 1bitaddie_1/inverter_1/out 1bitaddie_1/sum 0.20fF
C875 1bitaddie_2/ff_2/inverter_0/w_n8_n5# s2 0.03fF
C876 1bitaddie_1/ff_0/m1_58_n52# 1bitaddie_1/ff_0/m1_25_n37# 0.08fF
C877 1bitaddie_1/Bi 1bitaddie_1/xorg_0/pmos_1/w_n8_n5# 0.07fF
C878 1bitaddie_4/clk 1bitaddie_0/ff_2/m1_63_0# 0.27fF
C879 ff_1/nmos_3/a_0_n10# ff_1/inverter_0/in 0.05fF
C880 1bitaddie_0/sum 1bitaddie_0/xorg_1/m1_25_n11# 0.12fF
C881 1bitaddie_3/ff_1/pmos_2/w_n8_n5# vdd 0.08fF
C882 1bitaddie_3/inverter_0/out gnd 0.08fF
C883 1bitaddie_2/xorg_1/m1_102_n17# vdd 0.12fF
C884 1bitaddie_1/xorg_1/inverter_0/out 1bitaddie_1/xorg_1/A 0.25fF
C885 ff_1/m1_63_0# gnd 0.05fF
C886 1bitaddie_2/xorg_1/pmos_0/w_n8_n5# vdd 0.08fF
C887 ff_0/m1_106_n52# ff_0/inverter_0/in 0.08fF
C888 B4 1bitaddie_4/clk 0.17fF
C889 1bitaddie_4/ff_0/inverter_0/in 1bitaddie_4/clk 0.22fF
C890 1bitaddie_3/sum 1bitaddie_3/xorg_1/pmos_3/w_n8_n5# 0.03fF
C891 1bitaddie_2/inverter_1/out 1bitaddie_2/Cin 0.05fF
C892 1bitaddie_4/xorg_0/pmos_3/w_n8_n5# 1bitaddie_4/xorg_1/A 0.03fF
C893 1bitaddie_4/ff_2/m1_63_0# 1bitaddie_4/ff_2/m1_25_n37# 0.05fF
C894 1bitaddie_4/ff_2/m1_25_n37# gnd 0.08fF
C895 1bitaddie_4/ff_0/m1_58_n52# gnd 0.08fF
C896 1bitaddie_3/inverter_1/w_n8_n5# 1bitaddie_3/inverter_1/out 0.03fF
C897 gnd 1bitaddie_1/xorg_1/inverter_1/out 0.08fF
C898 1bitaddie_0/inverter_0/w_n8_n5# 1bitaddie_0/inverter_0/out 0.03fF
C899 1bitaddie_3/Ai 1bitaddie_3/ff_1/inverter_0/in 0.05fF
C900 1bitaddie_2/xorg_0/inverter_1/out 1bitaddie_2/xorg_0/m1_102_n91# 0.05fF
C901 1bitaddie_2/ff_2/inverter_0/in 1bitaddie_4/clk 0.05fF
C902 vdd 1bitaddie_1/inverter_1/w_n8_n5# 0.08fF
C903 1bitaddie_0/ff_0/m1_63_0# vdd 0.12fF
C904 1bitaddie_0/xorg_1/A inverter_0/out 0.10fF
C905 1bitaddie_1/manch_0/clk 1bitaddie_1/inverter_2/w_n8_n5# 0.03fF
C906 1bitaddie_0/ff_1/m1_58_n52# 1bitaddie_0/ff_1/m1_25_n37# 0.08fF
C907 1bitaddie_3/xorg_1/m1_102_n17# vdd 0.12fF
C908 1bitaddie_0/ff_2/inverter_0/in 1bitaddie_0/ff_2/pmos_3/w_n8_n5# 0.03fF
C909 A0 gnd 0.05fF
C910 1bitaddie_0/Ai 1bitaddie_0/xorg_0/m1_102_n17# 0.20fF
C911 1bitaddie_3/xorg_1/pmos_0/w_n8_n5# vdd 0.08fF
C912 1bitaddie_4/ff_1/inverter_0/w_n8_n5# vdd 0.08fF
C913 1bitaddie_0/sum 1bitaddie_0/ff_2/pmos_0/w_n8_n5# 0.07fF
C914 1bitaddie_4/sum 1bitaddie_4/clk 0.08fF
C915 ff_1/nmos_3/a_0_n10# ff_1/m1_106_n52# 0.05fF
C916 1bitaddie_1/inverter_1/out 1bitaddie_1/xorg_1/pmos_1/w_n8_n5# 0.07fF
C917 1bitaddie_0/ff_0/m1_25_n37# gnd 0.08fF
C918 1bitaddie_3/xorg_1/inverter_0/out 1bitaddie_3/xorg_1/A 0.25fF
C919 1bitaddie_2/ff_2/pmos_2/w_n8_n5# vdd 0.08fF
C920 1bitaddie_4/xorg_1/pmos_2/w_n8_n5# 1bitaddie_4/xorg_1/m1_102_n17# 0.03fF
C921 1bitaddie_3/ff_2/inverter_0/w_n8_n5# s3 0.03fF
C922 1bitaddie_3/ff_2/inverter_0/in 1bitaddie_4/clk 0.05fF
C923 1bitaddie_2/xorg_1/inverter_1/w_n8_n5# vdd 0.08fF
C924 1bitaddie_0/nandg_0/pmos_0/w_n8_n5# vdd 0.08fF
C925 1bitaddie_4/Ai 1bitaddie_4/Bi 0.06fF
C926 1bitaddie_4/ff_2/pmos_0/w_n8_n5# 1bitaddie_4/ff_2/m1_19_n10# 0.03fF
C927 1bitaddie_1/ff_1/pmos_3/w_n8_n5# 1bitaddie_1/ff_1/m1_63_0# 0.07fF
C928 1bitaddie_4/ff_2/inverter_0/in vdd 0.12fF
C929 B4 1bitaddie_4/ff_0/m1_25_n37# 0.05fF
C930 1bitaddie_4/Bi 1bitaddie_4/xorg_0/inverter_1/out 0.05fF
C931 1bitaddie_4/ff_1/inverter_0/w_n8_n5# 1bitaddie_4/ff_1/inverter_0/in 0.07fF
C932 m1_608_244# ff_0/m1_63_0# 0.05fF
C933 1bitaddie_3/inverter_1/out 1bitaddie_3/Cin 0.05fF
C934 1bitaddie_2/ff_0/inverter_0/w_n8_n5# 1bitaddie_2/ff_0/inverter_0/in 0.07fF
C935 1bitaddie_1/xorg_1/A 1bitaddie_1/xorg_1/m1_25_n11# 0.14fF
C936 1bitaddie_2/ff_2/m1_63_0# 1bitaddie_4/clk 0.27fF
C937 1bitaddie_1/xorg_0/pmos_1/w_n8_n5# 1bitaddie_1/xorg_0/m1_25_n11# 0.08fF
C938 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/xorg_1/m1_102_n91# 0.05fF
C939 1bitaddie_4/nandg_0/m1_26_n48# 1bitaddie_4/Ai 0.12fF
C940 1bitaddie_3/ff_2/pmos_2/w_n8_n5# vdd 0.08fF
C941 ff_1/inverter_0/in ff_1/m1_106_n52# 0.08fF
C942 1bitaddie_3/xorg_0/inverter_1/out 1bitaddie_3/xorg_0/m1_102_n91# 0.05fF
C943 1bitaddie_3/xorg_1/inverter_1/w_n8_n5# vdd 0.08fF
C944 1bitaddie_2/manch_0/m1_24_n50# 1bitaddie_2/manch_0/clk 0.05fF
C945 1bitaddie_2/xorg_0/m1_102_n91# 1bitaddie_2/xorg_1/A 0.08fF
C946 1bitaddie_0/ff_2/m1_63_0# 1bitaddie_0/ff_2/pmos_3/w_n8_n5# 0.07fF
C947 1bitaddie_1/manch_0/clk 1bitaddie_1/Cin 0.07fF
C948 1bitaddie_1/ff_1/inverter_0/w_n8_n5# 1bitaddie_1/ff_1/inverter_0/in 0.07fF
C949 vdd 1bitaddie_1/xorg_0/inverter_1/out 0.12fF
C950 1bitaddie_4/xorg_1/inverter_0/out gnd 0.14fF
C951 1bitaddie_0/nandg_0/m1_26_n48# 1bitaddie_0/Ai 0.12fF
C952 ff_1/pmos_1/w_n8_n5# ff_1/m1_19_n10# 0.08fF
C953 gnd 1bitaddie_1/ff_0/m1_63_0# 0.05fF
C954 1bitaddie_1/ff_1/m1_19_n10# A1 0.11fF
C955 1bitaddie_0/xorg_1/inverter_0/out 1bitaddie_0/xorg_1/pmos_0/w_n8_n5# 0.07fF
C956 1bitaddie_3/ff_2/m1_63_0# 1bitaddie_4/clk 0.27fF
C957 1bitaddie_2/ff_0/m1_63_0# vdd 0.12fF
C958 1bitaddie_1/xorg_0/m1_102_n91# 1bitaddie_1/xorg_1/A 0.08fF
C959 1bitaddie_2/manch_0/m1_24_n50# 1bitaddie_2/Cin 0.07fF
C960 1bitaddie_1/inverter_1/out 1bitaddie_1/inverter_1/w_n8_n5# 0.03fF
C961 1bitaddie_0/xorg_0/m1_102_n17# 1bitaddie_0/xorg_1/A 0.12fF
C962 1bitaddie_4/ff_2/m1_63_0# vdd 0.12fF
C963 1bitaddie_4/manch_0/pmos_0/w_n8_n5# inverter_1/out 0.03fF
C964 A2 gnd 0.05fF
C965 1bitaddie_2/ff_0/m1_63_0# 1bitaddie_2/ff_0/m1_25_n37# 0.05fF
C966 1bitaddie_1/Bi 1bitaddie_1/nandg_0/m1_26_n48# 0.05fF
C967 1bitaddie_0/ff_0/m1_63_0# 1bitaddie_0/ff_0/m1_58_n52# 0.08fF
C968 1bitaddie_4/xorg_0/inverter_0/out 1bitaddie_4/Ai 0.25fF
C969 1bitaddie_2/ff_0/m1_25_n37# gnd 0.08fF
C970 1bitaddie_0/ff_1/m1_25_n37# gnd 0.08fF
C971 1bitaddie_0/inverter_2/w_n8_n5# 1bitaddie_0/manch_0/clk 0.03fF
C972 1bitaddie_0/xorg_0/pmos_3/w_n8_n5# 1bitaddie_0/xorg_0/m1_102_n17# 0.08fF
C973 1bitaddie_3/ff_0/inverter_0/w_n8_n5# 1bitaddie_3/ff_0/inverter_0/in 0.07fF
C974 1bitaddie_0/ff_0/inverter_0/in 1bitaddie_0/ff_0/pmos_3/w_n8_n5# 0.03fF
C975 1bitaddie_4/Bi 1bitaddie_4/xorg_1/A 0.20fF
C976 1bitaddie_3/ff_0/m1_63_0# vdd 0.12fF
C977 1bitaddie_1/xorg_0/inverter_0/out 1bitaddie_1/xorg_1/A 0.06fF
C978 1bitaddie_4/clk 1bitaddie_1/ff_1/inverter_0/in 0.05fF
C979 1bitaddie_0/xorg_0/inverter_0/out 1bitaddie_0/xorg_0/m1_102_n91# 0.05fF
C980 1bitaddie_2/manch_0/m1_24_n50# 1bitaddie_3/Cin 0.08fF
C981 1bitaddie_4/Ai 1bitaddie_4/xorg_0/m1_25_n11# 0.14fF
C982 1bitaddie_4/sum 1bitaddie_4/ff_2/m1_19_n10# 0.11fF
C983 A3 gnd 0.05fF
C984 1bitaddie_3/manch_0/m1_24_n50# 1bitaddie_3/manch_0/clk 0.05fF
C985 1bitaddie_4/ff_1/inverter_0/in gnd 0.05fF
C986 1bitaddie_3/xorg_0/m1_102_n91# 1bitaddie_3/xorg_1/A 0.08fF
C987 1bitaddie_4/xorg_1/inverter_1/w_n8_n5# 1bitaddie_4/inverter_1/out 0.07fF
C988 inverter_1/w_n8_n5# inverter_1/out 0.03fF
C989 1bitaddie_4/clk 1bitaddie_1/ff_1/pmos_2/w_n8_n5# 0.07fF
C990 1bitaddie_0/xorg_1/pmos_1/w_n8_n5# 1bitaddie_0/xorg_1/m1_25_n11# 0.08fF
C991 1bitaddie_2/sum 1bitaddie_2/xorg_1/m1_25_n11# 0.12fF
C992 1bitaddie_3/ff_0/m1_25_n37# gnd 0.08fF
C993 1bitaddie_4/xorg_0/inverter_0/w_n8_n5# vdd 0.08fF
C994 1bitaddie_1/sum 1bitaddie_1/xorg_1/m1_102_n17# 0.12fF
C995 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/inverter_1/out 0.05fF
C996 1bitaddie_1/ff_1/pmos_1/w_n8_n5# 1bitaddie_1/ff_1/m1_19_n10# 0.08fF
C997 1bitaddie_3/manch_0/m1_24_n50# 1bitaddie_3/Cin 0.07fF
C998 1bitaddie_0/xorg_1/A 1bitaddie_0/xorg_1/pmos_2/w_n8_n5# 0.07fF
C999 1bitaddie_2/Bi 1bitaddie_2/nandg_0/pmos_0/w_n8_n5# 0.07fF
C1000 1bitaddie_4/ff_0/inverter_0/w_n8_n5# vdd 0.08fF
C1001 gnd 1bitaddie_1/ff_2/inverter_0/in 0.05fF
C1002 1bitaddie_3/ff_0/m1_63_0# 1bitaddie_3/ff_0/m1_25_n37# 0.05fF
C1003 1bitaddie_1/ff_0/m1_106_n52# 1bitaddie_1/ff_0/m1_63_0# 0.05fF
C1004 C0 ff_0/m1_19_n10# 0.11fF
C1005 1bitaddie_4/ff_2/inverter_0/in s4 0.05fF
C1006 1bitaddie_4/ff_1/pmos_0/w_n8_n5# vdd 0.08fF
C1007 1bitaddie_2/xorg_1/A 1bitaddie_2/Cin 0.10fF
C1008 1bitaddie_2/ff_1/m1_58_n52# 1bitaddie_2/ff_1/m1_25_n37# 0.08fF
C1009 1bitaddie_2/ff_2/inverter_0/in 1bitaddie_2/ff_2/pmos_3/w_n8_n5# 0.03fF
C1010 1bitaddie_2/Ai 1bitaddie_2/xorg_0/m1_102_n17# 0.20fF
C1011 1bitaddie_0/ff_2/m1_58_n52# 1bitaddie_0/ff_2/m1_25_n37# 0.08fF
C1012 1bitaddie_4/xorg_0/m1_102_n91# gnd 0.08fF
C1013 1bitaddie_4/inverter_0/in gnd 0.05fF
C1014 1bitaddie_2/sum 1bitaddie_2/ff_2/pmos_0/w_n8_n5# 0.07fF
C1015 1bitaddie_0/inverter_1/out 1bitaddie_0/xorg_1/m1_26_n95# 0.05fF
C1016 1bitaddie_4/xorg_1/inverter_0/out 1bitaddie_4/xorg_1/m1_25_n11# 0.05fF
C1017 gnd 1bitaddie_1/inverter_1/out 0.14fF
C1018 1bitaddie_4/clk B0 0.17fF
C1019 1bitaddie_4/clk 1bitaddie_0/ff_0/inverter_0/in 0.22fF
C1020 1bitaddie_4/xorg_0/inverter_0/out 1bitaddie_4/xorg_1/A 0.06fF
C1021 ff_1/pmos_1/w_n8_n5# ff_1/m1_25_n37# 0.03fF
C1022 1bitaddie_2/ff_1/m1_25_n37# gnd 0.08fF
C1023 gnd 1bitaddie_0/ff_2/m1_25_n37# 0.08fF
C1024 1bitaddie_0/ff_0/m1_58_n52# gnd 0.08fF
C1025 1bitaddie_1/ff_1/m1_25_n37# A1 0.05fF
C1026 1bitaddie_0/inverter_1/out 1bitaddie_0/xorg_1/A 0.06fF
C1027 1bitaddie_0/ff_1/m1_63_0# 1bitaddie_0/ff_1/pmos_2/w_n8_n5# 0.03fF
C1028 1bitaddie_3/sum 1bitaddie_3/xorg_1/m1_25_n11# 0.12fF
C1029 1bitaddie_2/xorg_1/A 1bitaddie_3/Cin 0.05fF
C1030 1bitaddie_4/xorg_0/m1_25_n11# 1bitaddie_4/xorg_1/A 0.12fF
C1031 1bitaddie_0/manch_0/clk 1bitaddie_1/Cin 0.16fF
C1032 1bitaddie_4/xorg_1/m1_25_n11# vdd 0.12fF
C1033 1bitaddie_1/xorg_0/inverter_0/w_n8_n5# vdd 0.08fF
C1034 vdd 1bitaddie_1/inverter_0/w_n8_n5# 0.08fF
C1035 1bitaddie_0/ff_1/inverter_0/w_n8_n5# vdd 0.08fF
C1036 1bitaddie_2/Ai 1bitaddie_2/nandg_0/pmos_1/w_n8_n5# 0.07fF
C1037 1bitaddie_0/ff_1/inverter_0/in 1bitaddie_0/ff_1/m1_106_n52# 0.08fF
C1038 1bitaddie_4/clk 1bitaddie_1/ff_2/pmos_2/w_n8_n5# 0.28fF
C1039 1bitaddie_1/ff_0/m1_19_n10# 1bitaddie_1/ff_0/m1_25_n37# 0.12fF
C1040 1bitaddie_4/clk 1bitaddie_0/sum 0.08fF
C1041 s4 gnd 0.08fF
C1042 gnd 1bitaddie_1/ff_2/m1_63_0# 0.05fF
C1043 B4 1bitaddie_4/ff_0/pmos_0/w_n8_n5# 0.07fF
C1044 1bitaddie_3/ff_1/m1_25_n37# gnd 0.08fF
C1045 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/xorg_1/m1_102_n91# 0.05fF
C1046 1bitaddie_2/Cin 1bitaddie_2/inverter_1/w_n8_n5# 0.07fF
C1047 inverter_0/out 1bitaddie_1/Cin 0.14fF
C1048 1bitaddie_0/inverter_0/w_n8_n5# vdd 0.08fF
C1049 1bitaddie_4/manch_0/pmos_0/w_n8_n5# vdd 0.08fF
C1050 1bitaddie_3/xorg_1/A 1bitaddie_3/Cin 0.10fF
C1051 1bitaddie_3/inverter_0/in 1bitaddie_3/inverter_0/w_n8_n5# 0.07fF
C1052 1bitaddie_2/ff_2/m1_63_0# 1bitaddie_2/ff_2/pmos_3/w_n8_n5# 0.07fF
C1053 1bitaddie_0/Bi 1bitaddie_0/xorg_0/m1_102_n17# 0.05fF
C1054 1bitaddie_4/ff_1/m1_63_0# gnd 0.05fF
C1055 1bitaddie_3/ff_1/m1_58_n52# 1bitaddie_3/ff_1/m1_25_n37# 0.08fF
C1056 1bitaddie_4/xorg_1/inverter_0/w_n8_n5# 1bitaddie_4/xorg_1/inverter_0/out 0.03fF
C1057 1bitaddie_3/ff_2/inverter_0/in 1bitaddie_3/ff_2/pmos_3/w_n8_n5# 0.03fF
C1058 1bitaddie_3/Ai 1bitaddie_3/xorg_0/m1_102_n17# 0.20fF
C1059 1bitaddie_0/ff_2/inverter_0/in vdd 0.12fF
C1060 1bitaddie_1/xorg_0/inverter_0/out 1bitaddie_1/Ai 0.25fF
C1061 1bitaddie_4/sum 1bitaddie_4/ff_2/m1_25_n37# 0.05fF
C1062 1bitaddie_2/xorg_1/inverter_0/out 1bitaddie_2/xorg_1/pmos_0/w_n8_n5# 0.07fF
C1063 1bitaddie_4/xorg_0/inverter_1/w_n8_n5# vdd 0.08fF
C1064 1bitaddie_3/sum 1bitaddie_3/ff_2/pmos_0/w_n8_n5# 0.07fF
C1065 ff_0/inverter_0/w_n8_n5# vdd 0.08fF
C1066 1bitaddie_4/ff_2/pmos_0/w_n8_n5# vdd 0.08fF
C1067 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/xorg_1/inverter_1/w_n8_n5# 0.03fF
C1068 1bitaddie_1/ff_1/inverter_0/in 1bitaddie_1/ff_1/m1_106_n52# 0.08fF
C1069 1bitaddie_4/xorg_1/A 1bitaddie_4/xorg_1/m1_102_n17# 0.20fF
C1070 1bitaddie_4/xorg_1/inverter_0/w_n8_n5# vdd 0.08fF
C1071 1bitaddie_4/manch_0/clk gnd 0.14fF
C1072 1bitaddie_2/xorg_0/m1_102_n17# 1bitaddie_2/xorg_1/A 0.12fF
C1073 1bitaddie_1/Cin 1bitaddie_1/xorg_1/A 0.10fF
C1074 1bitaddie_4/clk 1bitaddie_1/ff_0/pmos_2/w_n8_n5# 0.07fF
C1075 1bitaddie_1/ff_1/pmos_1/w_n8_n5# 1bitaddie_1/ff_1/m1_25_n37# 0.03fF
C1076 vdd 1bitaddie_1/xorg_1/pmos_0/w_n8_n5# 0.08fF
C1077 1bitaddie_0/ff_1/pmos_0/w_n8_n5# 1bitaddie_0/ff_1/m1_19_n10# 0.03fF
C1078 inverter_1/w_n8_n5# vdd 0.08fF
C1079 1bitaddie_2/ff_0/m1_63_0# 1bitaddie_2/ff_0/m1_58_n52# 0.08fF
C1080 1bitaddie_4/ff_0/m1_19_n10# 1bitaddie_4/clk 0.09fF
C1081 B2 1bitaddie_4/clk 0.17fF
C1082 1bitaddie_2/ff_0/inverter_0/in 1bitaddie_4/clk 0.22fF
C1083 1bitaddie_0/sum 1bitaddie_0/xorg_1/pmos_1/w_n8_n5# 0.03fF
C1084 1bitaddie_2/nandg_0/m1_26_n48# 1bitaddie_2/inverter_0/in 0.08fF
C1085 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_1/ff_2/m1_19_n10# 0.12fF
C1086 1bitaddie_0/xorg_1/inverter_0/out gnd 0.14fF
C1087 m1_641_206# C0 0.05fF
C1088 1bitaddie_2/ff_0/m1_58_n52# gnd 0.08fF
C1089 1bitaddie_2/xorg_0/pmos_3/w_n8_n5# 1bitaddie_2/xorg_0/m1_102_n17# 0.08fF
C1090 1bitaddie_2/ff_2/m1_25_n37# gnd 0.08fF
C1091 1bitaddie_1/xorg_0/m1_102_n17# 1bitaddie_1/xorg_1/A 0.12fF
C1092 1bitaddie_2/ff_0/inverter_0/in 1bitaddie_2/ff_0/pmos_3/w_n8_n5# 0.03fF
C1093 1bitaddie_1/xorg_1/inverter_0/out 1bitaddie_1/xorg_1/m1_102_n91# 0.05fF
C1094 1bitaddie_4/nandg_0/m1_26_n48# 1bitaddie_4/Bi 0.05fF
C1095 1bitaddie_4/Cin gnd 0.10fF
C1096 vdd 1bitaddie_1/Bi 0.24fF
C1097 1bitaddie_2/xorg_0/inverter_0/out 1bitaddie_2/xorg_0/m1_102_n91# 0.05fF
C1098 A0 1bitaddie_0/ff_1/pmos_0/w_n8_n5# 0.07fF
C1099 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/xorg_1/m1_102_n91# 0.05fF
C1100 vdd 1bitaddie_1/ff_2/inverter_0/w_n8_n5# 0.08fF
C1101 1bitaddie_3/ff_2/m1_63_0# 1bitaddie_3/ff_2/pmos_3/w_n8_n5# 0.07fF
C1102 1bitaddie_0/ff_2/m1_63_0# vdd 0.12fF
C1103 1bitaddie_0/inverter_0/in 1bitaddie_0/nandg_0/pmos_1/w_n8_n5# 0.03fF
C1104 1bitaddie_2/ff_1/inverter_0/w_n8_n5# vdd 0.08fF
C1105 1bitaddie_1/manch_0/pmos_0/w_n8_n5# vdd 0.08fF
C1106 1bitaddie_2/xorg_1/pmos_1/w_n8_n5# 1bitaddie_2/xorg_1/m1_25_n11# 0.08fF
C1107 1bitaddie_0/nandg_0/m1_26_n48# 1bitaddie_0/Bi 0.05fF
C1108 B3 1bitaddie_4/clk 0.17fF
C1109 1bitaddie_3/ff_0/inverter_0/in 1bitaddie_4/clk 0.22fF
C1110 1bitaddie_2/sum 1bitaddie_4/clk 0.08fF
C1111 1bitaddie_0/xorg_0/inverter_1/out 1bitaddie_0/xorg_1/A 0.22fF
C1112 1bitaddie_3/ff_0/m1_58_n52# gnd 0.08fF
C1113 1bitaddie_3/xorg_1/inverter_0/out 1bitaddie_3/xorg_1/pmos_0/w_n8_n5# 0.07fF
C1114 ff_1/m1_63_0# ff_1/pmos_2/w_n8_n5# 0.03fF
C1115 1bitaddie_3/ff_2/m1_25_n37# gnd 0.08fF
C1116 gnd 1bitaddie_1/xorg_0/m1_26_n95# 0.08fF
C1117 1bitaddie_2/Cin 1bitaddie_1/Cin 0.14fF
C1118 1bitaddie_2/xorg_1/inverter_1/out 1bitaddie_2/inverter_1/out 0.05fF
C1119 1bitaddie_0/xorg_0/inverter_0/out 1bitaddie_0/xorg_0/pmos_0/w_n8_n5# 0.07fF
C1120 1bitaddie_4/ff_0/inverter_0/in vdd 0.12fF
C1121 1bitaddie_1/xorg_0/inverter_1/w_n8_n5# vdd 0.08fF
C1122 1bitaddie_2/xorg_1/A 1bitaddie_2/xorg_1/pmos_2/w_n8_n5# 0.07fF
C1123 1bitaddie_1/ff_2/pmos_1/w_n8_n5# 1bitaddie_1/ff_2/m1_19_n10# 0.08fF
C1124 1bitaddie_4/ff_0/m1_19_n10# 1bitaddie_4/ff_0/m1_25_n37# 0.12fF
C1125 1bitaddie_3/xorg_0/m1_102_n17# 1bitaddie_3/xorg_1/A 0.12fF
C1126 1bitaddie_0/ff_1/m1_63_0# 1bitaddie_0/ff_1/m1_106_n52# 0.05fF
C1127 1bitaddie_0/xorg_0/inverter_1/out 1bitaddie_0/xorg_0/pmos_3/w_n8_n5# 0.07fF
C1128 1bitaddie_0/xorg_0/pmos_0/w_n8_n5# 1bitaddie_0/xorg_0/m1_25_n11# 0.03fF
C1129 1bitaddie_2/ff_2/inverter_0/in vdd 0.12fF
C1130 B0 1bitaddie_0/ff_0/m1_19_n10# 0.11fF
C1131 1bitaddie_1/manch_0/clk gnd 0.14fF
C1132 1bitaddie_3/ff_0/m1_63_0# 1bitaddie_3/ff_0/m1_58_n52# 0.08fF
C1133 1bitaddie_0/ff_1/inverter_0/in gnd 0.05fF
C1134 1bitaddie_3/ff_1/inverter_0/w_n8_n5# vdd 0.08fF
C1135 1bitaddie_3/Ai 1bitaddie_3/nandg_0/m1_26_n48# 0.12fF
C1136 1bitaddie_3/sum 1bitaddie_4/clk 0.08fF
C1137 1bitaddie_0/ff_1/m1_63_0# 1bitaddie_0/ff_1/m1_58_n52# 0.08fF
C1138 1bitaddie_3/xorg_0/pmos_3/w_n8_n5# 1bitaddie_3/xorg_0/m1_102_n17# 0.08fF
C1139 1bitaddie_1/xorg_1/inverter_0/out 1bitaddie_1/xorg_1/m1_25_n11# 0.05fF
C1140 1bitaddie_0/xorg_0/inverter_0/w_n8_n5# vdd 0.08fF
C1141 ff_1/nmos_3/a_0_n10# ff_1/m1_63_0# 0.02fF
C1142 1bitaddie_3/ff_0/inverter_0/in 1bitaddie_3/ff_0/pmos_3/w_n8_n5# 0.03fF
C1143 1bitaddie_4/clk 1bitaddie_1/ff_2/m1_106_n52# 0.05fF
C1144 1bitaddie_1/ff_2/inverter_0/in 1bitaddie_1/ff_2/inverter_0/w_n8_n5# 0.07fF
C1145 1bitaddie_2/ff_2/m1_58_n52# 1bitaddie_2/ff_2/m1_25_n37# 0.08fF
C1146 m1_560_235# ff_0/m1_63_0# 0.05fF
C1147 1bitaddie_3/xorg_0/inverter_0/out 1bitaddie_3/xorg_0/m1_102_n91# 0.05fF
C1148 1bitaddie_2/inverter_1/out 1bitaddie_2/xorg_1/m1_26_n95# 0.05fF
C1149 1bitaddie_4/ff_1/m1_19_n10# 1bitaddie_4/clk 0.09fF
C1150 1bitaddie_1/xorg_0/pmos_2/w_n8_n5# 1bitaddie_1/xorg_0/m1_102_n17# 0.03fF
C1151 1bitaddie_0/ff_0/inverter_0/w_n8_n5# vdd 0.08fF
C1152 1bitaddie_3/ff_2/inverter_0/in vdd 0.12fF
C1153 1bitaddie_2/manch_0/clk 1bitaddie_2/inverter_2/w_n8_n5# 0.03fF
C1154 1bitaddie_4/clk 1bitaddie_1/ff_2/m1_58_n52# 0.11fF
C1155 1bitaddie_2/xorg_1/inverter_0/out gnd 0.14fF
C1156 1bitaddie_3/xorg_1/pmos_1/w_n8_n5# 1bitaddie_3/xorg_1/m1_25_n11# 0.08fF
C1157 B1 1bitaddie_1/ff_0/m1_19_n10# 0.11fF
C1158 1bitaddie_0/xorg_1/m1_26_n95# 1bitaddie_0/xorg_1/A 0.05fF
C1159 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_2/ff_1/pmos_2/w_n8_n5# 0.03fF
C1160 1bitaddie_1/ff_1/m1_25_n37# 1bitaddie_1/ff_1/m1_63_0# 0.05fF
C1161 inverter_1/in gnd 0.11fF
C1162 1bitaddie_2/inverter_1/out 1bitaddie_2/xorg_1/A 0.06fF
C1163 1bitaddie_0/ff_1/pmos_0/w_n8_n5# vdd 0.08fF
C1164 vdd 1bitaddie_1/xorg_0/m1_25_n11# 0.12fF
C1165 A4 1bitaddie_4/clk 0.17fF
C1166 1bitaddie_1/xorg_1/inverter_1/out 1bitaddie_1/xorg_1/inverter_1/w_n8_n5# 0.03fF
C1167 1bitaddie_3/xorg_1/inverter_1/out 1bitaddie_3/inverter_1/out 0.05fF
C1168 1bitaddie_3/xorg_1/A 1bitaddie_3/xorg_1/pmos_2/w_n8_n5# 0.07fF
C1169 1bitaddie_2/ff_2/m1_63_0# vdd 0.12fF
C1170 ff_1/inverter_0/in ff_1/m1_63_0# 0.05fF
C1171 1bitaddie_0/xorg_0/m1_102_n91# gnd 0.08fF
C1172 1bitaddie_4/ff_0/pmos_3/w_n8_n5# vdd 0.06fF
C1173 1bitaddie_2/ff_1/inverter_0/in 1bitaddie_2/ff_1/m1_106_n52# 0.08fF
C1174 1bitaddie_4/ff_0/m1_25_n37# 1bitaddie_4/clk 0.31fF
C1175 1bitaddie_1/manch_0/m1_24_n50# 1bitaddie_1/Cin 0.07fF
C1176 1bitaddie_1/ff_0/pmos_0/w_n8_n5# 1bitaddie_1/ff_0/m1_19_n10# 0.03fF
C1177 1bitaddie_3/xorg_1/inverter_0/out gnd 0.14fF
C1178 1bitaddie_1/Bi 1bitaddie_1/ff_0/inverter_0/w_n8_n5# 0.03fF
C1179 A4 1bitaddie_4/ff_1/m1_19_n10# 0.11fF
C1180 1bitaddie_4/xorg_1/m1_102_n91# gnd 0.08fF
C1181 1bitaddie_0/xorg_0/pmos_3/w_n8_n5# 1bitaddie_0/xorg_1/A 0.03fF
C1182 1bitaddie_4/manch_0/pmos_0/w_n8_n5# 1bitaddie_4/manch_0/clk 0.07fF
C1183 1bitaddie_0/ff_2/m1_63_0# 1bitaddie_0/ff_2/m1_25_n37# 0.05fF
C1184 1bitaddie_0/inverter_0/in 1bitaddie_0/inverter_0/out 0.05fF
C1185 1bitaddie_2/Bi 1bitaddie_2/xorg_0/m1_102_n17# 0.05fF
C1186 1bitaddie_1/ff_0/pmos_1/w_n8_n5# 1bitaddie_1/ff_0/m1_19_n10# 0.08fF
C1187 1bitaddie_1/Ai 1bitaddie_1/xorg_0/m1_102_n17# 0.20fF
C1188 1bitaddie_3/ff_2/m1_58_n52# 1bitaddie_3/ff_2/m1_25_n37# 0.08fF
C1189 1bitaddie_0/xorg_1/m1_25_n11# vdd 0.12fF
C1190 1bitaddie_3/ff_2/m1_63_0# vdd 0.12fF
C1191 1bitaddie_4/inverter_0/out inverter_1/out 0.19fF
C1192 1bitaddie_3/inverter_1/out 1bitaddie_3/xorg_1/m1_26_n95# 0.05fF
C1193 1bitaddie_2/ff_1/inverter_0/in gnd 0.05fF
C1194 1bitaddie_3/inverter_0/w_n8_n5# 1bitaddie_3/inverter_0/out 0.03fF
C1195 1bitaddie_4/xorg_0/inverter_0/out 1bitaddie_4/xorg_0/m1_25_n11# 0.05fF
C1196 1bitaddie_2/inverter_1/out 1bitaddie_2/inverter_1/w_n8_n5# 0.03fF
C1197 s0 gnd 0.08fF
C1198 ff_1/pmos_2/w_n8_n5# vdd 0.08fF
C1199 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_3/ff_1/pmos_2/w_n8_n5# 0.03fF
C1200 1bitaddie_2/xorg_0/inverter_0/w_n8_n5# vdd 0.08fF
C1201 1bitaddie_3/inverter_1/out 1bitaddie_3/xorg_1/A 0.06fF
C1202 1bitaddie_0/xorg_1/pmos_2/w_n8_n5# 1bitaddie_0/xorg_1/m1_102_n17# 0.03fF
C1203 1bitaddie_0/manch_0/pmos_0/w_n8_n5# vdd 0.08fF
C1204 ff_1/m1_63_0# ff_1/m1_106_n52# 0.05fF
C1205 1bitaddie_2/ff_1/pmos_0/w_n8_n5# 1bitaddie_2/ff_1/m1_19_n10# 0.03fF
C1206 1bitaddie_0/Ai 1bitaddie_0/Bi 0.06fF
C1207 1bitaddie_0/ff_2/pmos_0/w_n8_n5# 1bitaddie_0/ff_2/m1_19_n10# 0.03fF
C1208 1bitaddie_0/ff_1/m1_63_0# gnd 0.05fF
C1209 1bitaddie_2/ff_0/inverter_0/w_n8_n5# vdd 0.08fF
C1210 1bitaddie_2/sum 1bitaddie_2/xorg_1/pmos_1/w_n8_n5# 0.03fF
C1211 vdd 1bitaddie_1/ff_1/inverter_0/in 0.12fF
C1212 1bitaddie_1/sum 1bitaddie_1/xorg_1/pmos_3/w_n8_n5# 0.03fF
C1213 B0 1bitaddie_0/ff_0/m1_25_n37# 0.05fF
C1214 C0 ff_0/m1_25_n37# 0.05fF
C1215 1bitaddie_3/ff_1/inverter_0/in 1bitaddie_3/ff_1/m1_106_n52# 0.08fF
C1216 1bitaddie_3/ff_1/inverter_0/in gnd 0.05fF
C1217 ff_1/m1_63_0# ff_1/m1_58_n52# 0.08fF
C1218 1bitaddie_0/Bi 1bitaddie_0/xorg_0/inverter_1/out 0.05fF
C1219 1bitaddie_0/xorg_0/inverter_1/w_n8_n5# vdd 0.08fF
C1220 1bitaddie_0/ff_1/inverter_0/w_n8_n5# 1bitaddie_0/ff_1/inverter_0/in 0.07fF
C1221 A2 1bitaddie_2/ff_1/pmos_0/w_n8_n5# 0.07fF
C1222 1bitaddie_2/ff_1/pmos_0/w_n8_n5# vdd 0.08fF
C1223 vdd 1bitaddie_0/ff_2/pmos_0/w_n8_n5# 0.08fF
C1224 1bitaddie_1/ff_2/m1_19_n10# 1bitaddie_1/sum 0.11fF
C1225 1bitaddie_1/Ai 1bitaddie_1/inverter_0/in 0.13fF
C1226 1bitaddie_3/xorg_0/inverter_0/w_n8_n5# vdd 0.08fF
C1227 1bitaddie_0/xorg_1/inverter_0/w_n8_n5# vdd 0.08fF
C1228 1bitaddie_4/ff_2/inverter_0/in 1bitaddie_4/ff_2/inverter_0/w_n8_n5# 0.07fF
C1229 vdd 1bitaddie_1/ff_1/pmos_2/w_n8_n5# 0.08fF
C1230 1bitaddie_0/manch_0/clk gnd 0.14fF
C1231 1bitaddie_3/Bi 1bitaddie_3/xorg_0/m1_102_n17# 0.05fF
C1232 1bitaddie_4/ff_1/pmos_3/w_n8_n5# vdd 0.06fF
C1233 1bitaddie_2/xorg_0/m1_102_n91# gnd 0.08fF
C1234 1bitaddie_4/clk 1bitaddie_0/ff_0/m1_19_n10# 0.09fF
C1235 1bitaddie_3/ff_0/inverter_0/w_n8_n5# vdd 0.08fF
C1236 gnd 1bitaddie_1/ff_0/m1_58_n52# 0.08fF
C1237 1bitaddie_4/ff_1/m1_25_n37# 1bitaddie_4/clk 0.41fF
C1238 1bitaddie_4/clk 1bitaddie_1/ff_1/m1_106_n52# 0.05fF
C1239 1bitaddie_2/xorg_0/inverter_1/out 1bitaddie_2/xorg_1/A 0.22fF
C1240 vdd 1bitaddie_1/xorg_1/inverter_1/w_n8_n5# 0.08fF
C1241 1bitaddie_4/inverter_1/out gnd 0.14fF
C1242 1bitaddie_2/xorg_0/inverter_0/out 1bitaddie_2/xorg_0/pmos_0/w_n8_n5# 0.07fF
C1243 B1 1bitaddie_1/ff_0/m1_25_n37# 0.05fF
C1244 gnd inverter_0/out 0.14fF
C1245 1bitaddie_3/ff_1/pmos_0/w_n8_n5# vdd 0.08fF
C1246 1bitaddie_4/clk 1bitaddie_1/ff_1/m1_58_n52# 0.12fF
C1247 ff_0/pmos_0/w_n8_n5# vdd 0.08fF
C1248 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_2/ff_1/m1_106_n52# 0.05fF
C1249 1bitaddie_2/xorg_0/inverter_1/out 1bitaddie_2/xorg_0/pmos_3/w_n8_n5# 0.07fF
C1250 1bitaddie_2/xorg_0/pmos_0/w_n8_n5# 1bitaddie_2/xorg_0/m1_25_n11# 0.03fF
C1251 1bitaddie_4/ff_1/m1_19_n10# 1bitaddie_4/ff_1/m1_25_n37# 0.12fF
C1252 B2 1bitaddie_2/ff_0/m1_19_n10# 0.11fF
C1253 1bitaddie_2/xorg_1/m1_25_n11# vdd 0.12fF
C1254 1bitaddie_1/xorg_0/inverter_1/out 1bitaddie_1/xorg_1/A 0.22fF
C1255 1bitaddie_4/Ai 1bitaddie_4/ff_1/inverter_0/w_n8_n5# 0.03fF
C1256 ff_1/inverter_0/in vdd 0.12fF
C1257 1bitaddie_3/ff_1/pmos_0/w_n8_n5# 1bitaddie_3/ff_1/m1_19_n10# 0.03fF
C1258 1bitaddie_1/Bi 1bitaddie_1/xorg_0/m1_26_n95# 0.05fF
C1259 1bitaddie_3/xorg_0/m1_102_n91# gnd 0.08fF
C1260 1bitaddie_2/inverter_0/out 1bitaddie_2/inverter_0/in 0.05fF
C1261 1bitaddie_4/ff_1/inverter_0/in 1bitaddie_4/ff_1/pmos_3/w_n8_n5# 0.03fF
C1262 1bitaddie_3/sum 1bitaddie_3/xorg_1/pmos_1/w_n8_n5# 0.03fF
C1263 gnd 1bitaddie_1/ff_0/inverter_0/in 0.05fF
C1264 1bitaddie_4/ff_0/pmos_1/w_n8_n5# 1bitaddie_4/ff_0/m1_19_n10# 0.08fF
C1265 1bitaddie_4/ff_0/pmos_0/w_n8_n5# 1bitaddie_4/ff_0/m1_19_n10# 0.03fF
C1266 1bitaddie_4/xorg_1/inverter_1/out 1bitaddie_4/xorg_1/pmos_3/w_n8_n5# 0.07fF
C1267 1bitaddie_4/xorg_0/pmos_1/w_n8_n5# 1bitaddie_4/xorg_1/A 0.03fF
C1268 1bitaddie_2/ff_1/m1_63_0# 1bitaddie_2/ff_1/m1_58_n52# 0.08fF
C1269 s2 gnd 0.08fF
C1270 m1_611_197# gnd 0.05fF
C1271 A4 1bitaddie_4/ff_1/m1_25_n37# 0.05fF
C1272 1bitaddie_1/xorg_0/inverter_0/out 1bitaddie_1/xorg_0/m1_102_n91# 0.05fF
C1273 1bitaddie_0/xorg_0/inverter_0/out 1bitaddie_0/Ai 0.25fF
C1274 1bitaddie_1/nandg_0/pmos_1/w_n8_n5# vdd 0.08fF
C1275 A3 1bitaddie_3/ff_1/pmos_0/w_n8_n5# 0.07fF
C1276 1bitaddie_0/ff_0/inverter_0/in vdd 0.12fF
C1277 1bitaddie_2/manch_0/pmos_0/w_n8_n5# vdd 0.08fF
C1278 gnd 1bitaddie_1/xorg_1/A 0.48fF
C1279 1bitaddie_0/Bi 1bitaddie_0/xorg_1/A 0.20fF
C1280 inverter_1/out 1bitaddie_4/clk 0.11fF
C1281 1bitaddie_4/ff_0/m1_63_0# 1bitaddie_4/ff_0/pmos_2/w_n8_n5# 0.03fF
C1282 1bitaddie_2/ff_1/m1_63_0# gnd 0.05fF
C1283 1bitaddie_1/ff_0/pmos_1/w_n8_n5# 1bitaddie_1/ff_0/m1_25_n37# 0.03fF
C1284 1bitaddie_0/Ai 1bitaddie_0/xorg_0/m1_25_n11# 0.14fF
C1285 1bitaddie_0/manch_0/m1_24_n50# 1bitaddie_1/Cin 0.08fF
C1286 1bitaddie_3/xorg_1/m1_25_n11# vdd 0.12fF
C1287 1bitaddie_1/manch_0/pmos_0/w_n8_n5# 1bitaddie_1/manch_0/clk 0.07fF
C1288 1bitaddie_2/xorg_1/m1_26_n95# 1bitaddie_2/xorg_1/A 0.05fF
C1289 1bitaddie_0/sum 1bitaddie_0/ff_2/m1_19_n10# 0.11fF
C1290 1bitaddie_2/xorg_0/inverter_1/w_n8_n5# vdd 0.08fF
C1291 1bitaddie_0/xorg_1/inverter_1/w_n8_n5# 1bitaddie_0/inverter_1/out 0.07fF
C1292 1bitaddie_3/xorg_0/inverter_1/out 1bitaddie_3/xorg_1/A 0.22fF
C1293 inverter_1/w_n8_n5# inverter_1/in 0.07fF
C1294 1bitaddie_3/inverter_0/w_n8_n5# vdd 0.08fF
C1295 s3 gnd 0.08fF
C1296 1bitaddie_3/inverter_2/w_n8_n5# 1bitaddie_4/clk 0.07fF
C1297 1bitaddie_2/ff_2/pmos_0/w_n8_n5# vdd 0.08fF
C1298 1bitaddie_3/xorg_0/inverter_0/out 1bitaddie_3/xorg_0/pmos_0/w_n8_n5# 0.07fF
C1299 1bitaddie_2/xorg_1/inverter_0/w_n8_n5# vdd 0.08fF
C1300 1bitaddie_2/manch_0/clk gnd 0.14fF
C1301 vdd 1bitaddie_1/ff_2/pmos_2/w_n8_n5# 0.08fF
C1302 1bitaddie_4/inverter_0/out vdd 0.12fF
C1303 1bitaddie_3/manch_0/pmos_0/w_n8_n5# vdd 0.08fF
C1304 1bitaddie_4/ff_2/pmos_3/w_n8_n5# vdd 0.06fF
C1305 1bitaddie_3/ff_1/m1_63_0# gnd 0.05fF
C1306 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_3/ff_1/m1_106_n52# 0.05fF
C1307 1bitaddie_2/ff_0/m1_19_n10# 1bitaddie_4/clk 0.09fF
C1308 1bitaddie_4/clk 1bitaddie_0/ff_1/m1_19_n10# 0.09fF
C1309 B3 1bitaddie_3/ff_0/m1_19_n10# 0.11fF
C1310 1bitaddie_3/xorg_0/inverter_1/out 1bitaddie_3/xorg_0/pmos_3/w_n8_n5# 0.07fF
C1311 1bitaddie_3/xorg_0/pmos_0/w_n8_n5# 1bitaddie_3/xorg_0/m1_25_n11# 0.03fF
C1312 1bitaddie_4/clk 1bitaddie_4/ff_2/m1_25_n37# 0.27fF
C1313 1bitaddie_4/ff_0/m1_58_n52# 1bitaddie_4/clk 0.12fF
C1314 1bitaddie_3/Bi 1bitaddie_3/nandg_0/m1_26_n48# 0.05fF
C1315 1bitaddie_3/inverter_0/in 1bitaddie_3/inverter_0/out 0.05fF
C1316 1bitaddie_2/xorg_0/pmos_3/w_n8_n5# 1bitaddie_2/xorg_1/A 0.03fF
C1317 1bitaddie_2/ff_2/m1_63_0# 1bitaddie_2/ff_2/m1_25_n37# 0.05fF
C1318 1bitaddie_3/xorg_0/inverter_1/w_n8_n5# vdd 0.08fF
C1319 1bitaddie_3/ff_1/m1_63_0# 1bitaddie_3/ff_1/m1_58_n52# 0.08fF
C1320 1bitaddie_2/Cin gnd 0.10fF
C1321 1bitaddie_1/xorg_1/inverter_1/w_n8_n5# 1bitaddie_1/inverter_1/out 0.07fF
C1322 1bitaddie_4/ff_0/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.30fF
C1323 inverter_0/w_n8_n5# vdd 0.08fF
C1324 1bitaddie_1/ff_0/m1_63_0# 1bitaddie_1/ff_0/pmos_2/w_n8_n5# 0.03fF
C1325 1bitaddie_0/ff_2/inverter_0/in s0 0.05fF
C1326 1bitaddie_3/ff_2/pmos_0/w_n8_n5# vdd 0.08fF
C1327 ff_0/inverter_0/in vdd 0.12fF
C1328 1bitaddie_4/clk A0 0.17fF
C1329 1bitaddie_4/Ai gnd 0.27fF
C1330 1bitaddie_3/xorg_1/inverter_0/w_n8_n5# vdd 0.08fF
C1331 1bitaddie_3/manch_0/clk gnd 0.14fF
C1332 1bitaddie_4/manch_0/m1_24_n50# gnd 0.08fF
C1333 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_1/ff_2/pmos_1/w_n8_n5# 0.03fF
C1334 1bitaddie_1/xorg_0/pmos_3/w_n8_n5# 1bitaddie_1/xorg_1/A 0.03fF
C1335 1bitaddie_0/ff_0/pmos_3/w_n8_n5# vdd 0.06fF
C1336 1bitaddie_3/ff_0/m1_19_n10# 1bitaddie_4/clk 0.09fF
C1337 1bitaddie_1/ff_0/m1_106_n52# 1bitaddie_1/ff_0/inverter_0/in 0.08fF
C1338 1bitaddie_4/clk 1bitaddie_0/ff_0/m1_25_n37# 0.31fF
C1339 1bitaddie_4/xorg_0/inverter_1/out gnd 0.08fF
C1340 vdd 1bitaddie_1/ff_0/pmos_2/w_n8_n5# 0.08fF
C1341 1bitaddie_0/xorg_1/inverter_0/out 1bitaddie_0/xorg_1/m1_25_n11# 0.05fF
C1342 ff_0/m1_25_n37# gnd 0.08fF
C1343 1bitaddie_3/xorg_1/m1_26_n95# 1bitaddie_3/xorg_1/A 0.05fF
C1344 1bitaddie_0/xorg_1/m1_102_n91# gnd 0.08fF
C1345 1bitaddie_4/ff_0/m1_19_n10# vdd 0.12fF
C1346 1bitaddie_1/sum 1bitaddie_1/xorg_1/m1_102_n91# 0.08fF
C1347 1bitaddie_0/xorg_0/inverter_0/out 1bitaddie_0/xorg_1/A 0.06fF
C1348 ff_1/nmos_2/a_0_n10# gnd 0.05fF
C1349 1bitaddie_3/Cin gnd 0.10fF
C1350 1bitaddie_2/xorg_1/pmos_2/w_n8_n5# 1bitaddie_2/xorg_1/m1_102_n17# 0.03fF
C1351 1bitaddie_2/ff_0/inverter_0/in vdd 0.12fF
C1352 1bitaddie_2/Ai 1bitaddie_2/Bi 0.06fF
C1353 1bitaddie_2/ff_2/pmos_0/w_n8_n5# 1bitaddie_2/ff_2/m1_19_n10# 0.03fF
C1354 1bitaddie_0/xorg_1/A 1bitaddie_1/Cin 0.05fF
C1355 1bitaddie_4/xorg_1/inverter_1/out gnd 0.08fF
C1356 1bitaddie_0/xorg_0/m1_25_n11# 1bitaddie_0/xorg_1/A 0.12fF
C1357 1bitaddie_4/ff_1/m1_63_0# 1bitaddie_4/ff_1/pmos_3/w_n8_n5# 0.07fF
C1358 1bitaddie_4/ff_0/m1_58_n52# 1bitaddie_4/ff_0/m1_25_n37# 0.08fF
C1359 B2 1bitaddie_2/ff_0/m1_25_n37# 0.05fF
C1360 1bitaddie_1/ff_1/inverter_0/w_n8_n5# vdd 0.08fF
C1361 1bitaddie_2/Bi 1bitaddie_2/xorg_0/inverter_1/out 0.05fF
C1362 1bitaddie_1/inverter_0/out vdd 0.12fF
C1363 1bitaddie_2/ff_1/inverter_0/w_n8_n5# 1bitaddie_2/ff_1/inverter_0/in 0.07fF
C1364 1bitaddie_4/ff_0/pmos_1/w_n8_n5# 1bitaddie_4/ff_0/m1_25_n37# 0.03fF
C1365 1bitaddie_4/xorg_0/inverter_0/w_n8_n5# 1bitaddie_4/Ai 0.07fF
C1366 1bitaddie_3/xorg_0/pmos_3/w_n8_n5# 1bitaddie_3/xorg_1/A 0.03fF
C1367 1bitaddie_3/ff_2/m1_63_0# 1bitaddie_3/ff_2/m1_25_n37# 0.05fF
C1368 B0 1bitaddie_0/ff_0/pmos_0/w_n8_n5# 0.07fF
C1369 1bitaddie_3/ff_0/inverter_0/in vdd 0.12fF
C1370 1bitaddie_0/inverter_0/in vdd 0.25fF
C1371 1bitaddie_4/inverter_0/in 1bitaddie_4/inverter_0/out 0.05fF
C1372 1bitaddie_2/ff_1/m1_19_n10# 1bitaddie_4/clk 0.09fF
C1373 1bitaddie_4/clk 1bitaddie_1/ff_0/m1_63_0# 0.35fF
C1374 1bitaddie_0/xorg_1/inverter_0/w_n8_n5# 1bitaddie_0/xorg_1/inverter_0/out 0.03fF
C1375 1bitaddie_0/nandg_0/m1_26_n48# gnd 0.08fF
C1376 1bitaddie_1/Ai gnd 0.27fF
C1377 1bitaddie_4/xorg_1/m1_102_n91# 1bitaddie_4/sum 0.08fF
C1378 1bitaddie_4/xorg_1/m1_26_n95# gnd 0.08fF
C1379 1bitaddie_1/manch_0/m1_24_n50# gnd 0.08fF
C1380 1bitaddie_4/Bi 1bitaddie_4/xorg_0/pmos_1/w_n8_n5# 0.07fF
C1381 1bitaddie_0/sum 1bitaddie_0/ff_2/m1_25_n37# 0.05fF
C1382 1bitaddie_0/nandg_0/pmos_1/w_n8_n5# vdd 0.08fF
C1383 B1 1bitaddie_1/ff_0/pmos_0/w_n8_n5# 0.07fF
C1384 vdd 1bitaddie_2/inverter_0/in 0.25fF
C1385 1bitaddie_1/sum 1bitaddie_1/xorg_1/m1_25_n11# 0.12fF
C1386 1bitaddie_4/ff_1/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.31fF
C1387 1bitaddie_0/xorg_1/inverter_1/out 1bitaddie_0/xorg_1/inverter_1/w_n8_n5# 0.03fF
C1388 1bitaddie_4/xorg_1/A gnd 0.48fF
C1389 A2 1bitaddie_4/clk 0.17fF
C1390 1bitaddie_4/clk vdd 0.43fF
C1391 1bitaddie_0/xorg_1/A 1bitaddie_0/xorg_1/m1_102_n17# 0.20fF
C1392 1bitaddie_4/ff_2/m1_19_n10# 1bitaddie_4/ff_2/m1_25_n37# 0.12fF
C1393 1bitaddie_3/xorg_1/pmos_2/w_n8_n5# 1bitaddie_3/xorg_1/m1_102_n17# 0.03fF
C1394 1bitaddie_4/ff_0/m1_106_n52# 1bitaddie_4/ff_0/m1_63_0# 0.05fF
C1395 1bitaddie_3/Ai 1bitaddie_3/Bi 0.06fF
C1396 1bitaddie_3/ff_2/pmos_0/w_n8_n5# 1bitaddie_3/ff_2/m1_19_n10# 0.03fF
C1397 1bitaddie_2/ff_0/pmos_3/w_n8_n5# vdd 0.06fF
C1398 1bitaddie_0/ff_1/pmos_3/w_n8_n5# vdd 0.06fF
C1399 1bitaddie_3/ff_1/m1_19_n10# 1bitaddie_4/clk 0.09fF
C1400 B3 1bitaddie_3/ff_0/m1_25_n37# 0.05fF
C1401 1bitaddie_2/ff_0/m1_25_n37# 1bitaddie_4/clk 0.31fF
C1402 1bitaddie_4/clk 1bitaddie_0/ff_1/m1_25_n37# 0.41fF
C1403 1bitaddie_1/ff_2/pmos_2/w_n8_n5# 1bitaddie_1/ff_2/m1_63_0# 0.03fF
C1404 1bitaddie_4/ff_1/pmos_1/w_n8_n5# 1bitaddie_4/ff_1/m1_19_n10# 0.08fF
C1405 ff_1/m1_25_n37# gnd 0.08fF
C1406 1bitaddie_3/Bi 1bitaddie_3/xorg_0/inverter_1/out 0.05fF
C1407 1bitaddie_2/xorg_1/m1_102_n91# gnd 0.08fF
C1408 1bitaddie_2/xorg_0/inverter_0/out 1bitaddie_2/Ai 0.25fF
C1409 1bitaddie_4/ff_1/m1_19_n10# vdd 0.12fF
C1410 1bitaddie_3/ff_1/inverter_0/w_n8_n5# 1bitaddie_3/ff_1/inverter_0/in 0.07fF
C1411 1bitaddie_0/inverter_1/out gnd 0.14fF
C1412 1bitaddie_3/inverter_0/in vdd 0.25fF
C1413 1bitaddie_2/Bi 1bitaddie_2/xorg_1/A 0.20fF
C1414 ff_0/m1_63_0# gnd 0.05fF
C1415 A3 1bitaddie_4/clk 0.17fF
C1416 1bitaddie_2/Ai 1bitaddie_2/xorg_0/m1_25_n11# 0.14fF
C1417 1bitaddie_1/Bi 1bitaddie_1/ff_0/inverter_0/in 0.05fF
C1418 1bitaddie_4/ff_1/inverter_0/in 1bitaddie_4/clk 0.05fF
C1419 1bitaddie_2/sum 1bitaddie_2/ff_2/m1_19_n10# 0.11fF
C1420 1bitaddie_3/ff_0/pmos_3/w_n8_n5# vdd 0.06fF
C1421 ff_0/pmos_0/w_n8_n5# ff_0/m1_19_n10# 0.03fF
C1422 1bitaddie_2/xorg_1/inverter_1/w_n8_n5# 1bitaddie_2/inverter_1/out 0.07fF
C1423 1bitaddie_3/ff_0/m1_25_n37# 1bitaddie_4/clk 0.31fF
C1424 1bitaddie_1/Bi 1bitaddie_1/xorg_1/A 0.20fF
C1425 1bitaddie_1/xorg_0/inverter_0/out 1bitaddie_1/xorg_0/pmos_0/w_n8_n5# 0.07fF
C1426 1bitaddie_3/xorg_1/m1_102_n91# gnd 0.08fF
C1427 gnd 1bitaddie_1/ff_1/m1_25_n37# 0.08fF
C1428 1bitaddie_1/xorg_1/pmos_1/w_n8_n5# 1bitaddie_1/xorg_1/m1_25_n11# 0.08fF
C1429 1bitaddie_4/inverter_0/out 1bitaddie_4/manch_0/clk 0.03fF
C1430 1bitaddie_1/ff_2/m1_25_n37# 1bitaddie_1/sum 0.05fF
C1431 1bitaddie_4/clk 1bitaddie_1/ff_2/inverter_0/in 0.05fF
C1432 1bitaddie_0/ff_0/m1_19_n10# 1bitaddie_0/ff_0/m1_25_n37# 0.12fF
C1433 1bitaddie_1/ff_2/m1_106_n52# 1bitaddie_1/ff_2/inverter_0/in 0.08fF
C1434 1bitaddie_1/ff_1/pmos_3/w_n8_n5# 1bitaddie_1/ff_1/inverter_0/in 0.03fF
C1435 1bitaddie_4/inverter_1/out 1bitaddie_4/sum 0.20fF
C1436 1bitaddie_4/xorg_0/pmos_1/w_n8_n5# 1bitaddie_4/xorg_0/m1_25_n11# 0.08fF
C1437 1bitaddie_3/manch_0/pmos_0/w_n8_n5# 1bitaddie_4/Cin 0.03fF
C1438 1bitaddie_1/xorg_1/m1_26_n95# 1bitaddie_1/inverter_1/out 0.05fF
C1439 1bitaddie_4/inverter_0/out 1bitaddie_4/Cin 0.02fF
C1440 1bitaddie_2/ff_2/inverter_0/in s2 0.05fF
C1441 ff_0/inverter_0/in ff_0/pmos_3/w_n8_n5# 0.03fF
C1442 1bitaddie_4/ff_2/pmos_1/w_n8_n5# 1bitaddie_4/clk 0.07fF
C1443 1bitaddie_4/xorg_0/inverter_1/w_n8_n5# 1bitaddie_4/xorg_0/inverter_1/out 0.03fF
C1444 1bitaddie_3/xorg_0/inverter_0/out 1bitaddie_3/Ai 0.25fF
C1445 vdd 1bitaddie_1/xorg_1/pmos_2/w_n8_n5# 0.08fF
C1446 ff_1/inverter_0/in ff_1/pmos_3/w_n8_n5# 0.03fF
C1447 1bitaddie_3/Bi 1bitaddie_3/xorg_1/A 0.20fF
C1448 1bitaddie_0/inverter_0/out vdd 0.12fF
C1449 1bitaddie_4/clk 1bitaddie_1/inverter_1/out 0.06fF
C1450 1bitaddie_4/xorg_0/pmos_2/w_n8_n5# vdd 0.08fF
C1451 1bitaddie_3/Ai 1bitaddie_3/xorg_0/m1_25_n11# 0.14fF
C1452 1bitaddie_2/ff_1/pmos_3/w_n8_n5# vdd 0.06fF
C1453 1bitaddie_1/xorg_0/inverter_0/w_n8_n5# 1bitaddie_1/Ai 0.07fF
C1454 vdd 1bitaddie_0/ff_2/pmos_3/w_n8_n5# 0.06fF
C1455 1bitaddie_2/ff_1/m1_25_n37# 1bitaddie_4/clk 0.41fF
C1456 1bitaddie_2/xorg_1/inverter_0/out 1bitaddie_2/xorg_1/m1_25_n11# 0.05fF
C1457 1bitaddie_4/clk 1bitaddie_0/ff_2/m1_25_n37# 0.27fF
C1458 1bitaddie_4/clk 1bitaddie_0/ff_0/m1_58_n52# 0.12fF
C1459 1bitaddie_3/sum 1bitaddie_3/ff_2/m1_19_n10# 0.11fF
C1460 1bitaddie_2/xorg_0/inverter_0/out 1bitaddie_2/xorg_1/A 0.06fF
C1461 1bitaddie_1/nandg_0/pmos_0/w_n8_n5# 1bitaddie_1/inverter_0/in 0.03fF
C1462 1bitaddie_3/xorg_1/inverter_1/w_n8_n5# 1bitaddie_3/inverter_1/out 0.07fF
C1463 1bitaddie_4/ff_2/m1_19_n10# vdd 0.12fF
C1464 1bitaddie_2/inverter_1/out gnd 0.14fF
C1465 1bitaddie_4/xorg_1/A 1bitaddie_4/xorg_1/m1_25_n11# 0.14fF
C1466 1bitaddie_1/manch_0/pmos_0/w_n8_n5# 1bitaddie_2/Cin 0.03fF
C1467 inverter_0/out Gnd 1.72fF
C1468 1bitaddie_0/ff_2/m1_25_n37# Gnd 0.41fF
C1469 1bitaddie_0/ff_2/pmos_3/w_n8_n5# Gnd 0.58fF
C1470 1bitaddie_0/ff_2/pmos_2/w_n8_n5# Gnd 0.58fF
C1471 1bitaddie_0/ff_2/m1_19_n10# Gnd 0.14fF
C1472 1bitaddie_0/ff_2/pmos_1/w_n8_n5# Gnd 0.58fF
C1473 1bitaddie_0/ff_2/pmos_0/w_n8_n5# Gnd 0.58fF
C1474 1bitaddie_0/ff_2/inverter_0/in Gnd 0.38fF
C1475 1bitaddie_0/ff_2/m1_106_n52# Gnd 0.26fF
C1476 1bitaddie_0/ff_2/m1_63_0# Gnd 0.69fF
C1477 1bitaddie_0/ff_2/m1_58_n52# Gnd 0.24fF
C1478 1bitaddie_0/ff_2/inverter_0/w_n8_n5# Gnd 0.53fF
C1479 gnd Gnd 23.71fF
C1480 1bitaddie_0/ff_1/m1_25_n37# Gnd 0.41fF
C1481 vdd Gnd 9.26fF
C1482 1bitaddie_0/ff_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1483 1bitaddie_0/ff_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1484 1bitaddie_0/ff_1/m1_19_n10# Gnd 0.14fF
C1485 1bitaddie_0/ff_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1486 1bitaddie_0/ff_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1487 1bitaddie_0/ff_1/inverter_0/in Gnd 0.38fF
C1488 1bitaddie_0/ff_1/m1_106_n52# Gnd 0.26fF
C1489 1bitaddie_0/ff_1/m1_63_0# Gnd 0.69fF
C1490 1bitaddie_0/ff_1/m1_58_n52# Gnd 0.24fF
C1491 A0 Gnd 0.54fF
C1492 1bitaddie_0/ff_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1493 1bitaddie_0/ff_0/m1_25_n37# Gnd 0.41fF
C1494 1bitaddie_0/ff_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1495 1bitaddie_0/ff_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1496 1bitaddie_0/ff_0/m1_19_n10# Gnd 0.14fF
C1497 1bitaddie_0/ff_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1498 1bitaddie_0/ff_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1499 1bitaddie_0/ff_0/inverter_0/in Gnd 0.38fF
C1500 1bitaddie_0/ff_0/m1_106_n52# Gnd 0.26fF
C1501 1bitaddie_0/ff_0/m1_63_0# Gnd 0.69fF
C1502 1bitaddie_0/ff_0/m1_58_n52# Gnd 0.24fF
C1503 B0 Gnd 0.59fF
C1504 1bitaddie_0/ff_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1505 1bitaddie_0/xorg_1/m1_102_n17# Gnd 0.04fF
C1506 1bitaddie_0/xorg_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1507 1bitaddie_0/xorg_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1508 1bitaddie_0/xorg_1/m1_25_n11# Gnd 0.13fF
C1509 1bitaddie_0/xorg_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1510 1bitaddie_0/xorg_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1511 1bitaddie_0/xorg_1/m1_102_n91# Gnd 0.22fF
C1512 1bitaddie_0/xorg_1/inverter_1/out Gnd 0.45fF
C1513 1bitaddie_0/sum Gnd 1.47fF
C1514 1bitaddie_0/xorg_1/m1_26_n95# Gnd 0.22fF
C1515 1bitaddie_0/inverter_1/out Gnd 0.90fF
C1516 1bitaddie_0/xorg_1/inverter_1/w_n8_n5# Gnd 0.53fF
C1517 1bitaddie_0/xorg_1/inverter_0/out Gnd 1.68fF
C1518 1bitaddie_0/xorg_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1519 1bitaddie_0/xorg_0/m1_102_n17# Gnd 0.04fF
C1520 1bitaddie_0/xorg_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1521 1bitaddie_0/xorg_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1522 1bitaddie_0/xorg_0/m1_25_n11# Gnd 0.13fF
C1523 1bitaddie_0/xorg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1524 1bitaddie_0/xorg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1525 1bitaddie_0/xorg_0/m1_102_n91# Gnd 0.22fF
C1526 1bitaddie_0/xorg_0/inverter_1/out Gnd 0.45fF
C1527 1bitaddie_0/xorg_0/m1_26_n95# Gnd 0.22fF
C1528 1bitaddie_0/Bi Gnd 1.53fF
C1529 1bitaddie_0/xorg_0/inverter_1/w_n8_n5# Gnd 0.53fF
C1530 1bitaddie_0/xorg_0/inverter_0/out Gnd 1.68fF
C1531 1bitaddie_0/Ai Gnd 2.80fF
C1532 1bitaddie_0/xorg_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1533 1bitaddie_0/manch_0/clk Gnd 1.66fF
C1534 1bitaddie_0/manch_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1535 1bitaddie_0/manch_0/m1_24_n50# Gnd 0.22fF
C1536 1bitaddie_0/inverter_0/out Gnd 0.59fF
C1537 1bitaddie_0/inverter_2/w_n8_n5# Gnd 0.53fF
C1538 1bitaddie_0/inverter_1/w_n8_n5# Gnd 0.53fF
C1539 1bitaddie_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1540 1bitaddie_0/inverter_0/in Gnd 1.07fF
C1541 1bitaddie_0/nandg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1542 1bitaddie_0/nandg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1543 1bitaddie_0/nandg_0/m1_26_n48# Gnd 0.21fF
C1544 ff_1/m1_25_n37# Gnd 0.41fF
C1545 ff_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1546 ff_1/pmos_2/a_0_n10# Gnd 0.11fF
C1547 ff_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1548 ff_1/m1_19_n10# Gnd 0.14fF
C1549 ff_1/pmos_1/a_0_n10# Gnd 0.11fF
C1550 ff_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1551 ff_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1552 ff_1/inverter_0/in Gnd 0.38fF
C1553 ff_1/m1_106_n52# Gnd 0.26fF
C1554 ff_1/nmos_3/a_0_n10# Gnd 0.16fF
C1555 ff_1/nmos_2/a_0_n10# Gnd 0.16fF
C1556 ff_1/m1_63_0# Gnd 0.69fF
C1557 ff_1/m1_58_n52# Gnd 0.24fF
C1558 inverter_1/in Gnd 0.77fF
C1559 Cout Gnd 0.11fF
C1560 ff_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1561 ff_0/m1_25_n37# Gnd 0.41fF
C1562 ff_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1563 m1_608_244# Gnd 0.17fF
C1564 ff_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1565 ff_0/m1_19_n10# Gnd 0.14fF
C1566 m1_641_206# Gnd 0.10fF
C1567 ff_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1568 ff_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1569 ff_0/inverter_0/in Gnd 0.38fF
C1570 ff_0/m1_106_n52# Gnd 0.26fF
C1571 m1_560_235# Gnd 0.29fF
C1572 ff_0/m1_63_0# Gnd 0.69fF
C1573 ff_0/m1_58_n52# Gnd 0.24fF
C1574 C0 Gnd 0.54fF
C1575 ff_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1576 1bitaddie_4/Cin Gnd 4.41fF
C1577 1bitaddie_4/ff_2/m1_25_n37# Gnd 0.41fF
C1578 1bitaddie_4/ff_2/pmos_3/w_n8_n5# Gnd 0.58fF
C1579 1bitaddie_4/clk Gnd 17.50fF
C1580 1bitaddie_4/ff_2/pmos_2/w_n8_n5# Gnd 0.58fF
C1581 1bitaddie_4/ff_2/m1_19_n10# Gnd 0.14fF
C1582 1bitaddie_4/ff_2/pmos_1/w_n8_n5# Gnd 0.58fF
C1583 1bitaddie_4/ff_2/pmos_0/w_n8_n5# Gnd 0.58fF
C1584 1bitaddie_4/ff_2/inverter_0/in Gnd 0.38fF
C1585 1bitaddie_4/ff_2/m1_106_n52# Gnd 0.26fF
C1586 1bitaddie_4/ff_2/m1_63_0# Gnd 0.69fF
C1587 1bitaddie_4/ff_2/m1_58_n52# Gnd 0.24fF
C1588 1bitaddie_4/ff_2/inverter_0/w_n8_n5# Gnd 0.53fF
C1589 1bitaddie_4/ff_1/m1_25_n37# Gnd 0.41fF
C1590 1bitaddie_4/ff_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1591 1bitaddie_4/ff_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1592 1bitaddie_4/ff_1/m1_19_n10# Gnd 0.14fF
C1593 1bitaddie_4/ff_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1594 1bitaddie_4/ff_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1595 1bitaddie_4/ff_1/inverter_0/in Gnd 0.38fF
C1596 1bitaddie_4/ff_1/m1_106_n52# Gnd 0.26fF
C1597 1bitaddie_4/ff_1/m1_63_0# Gnd 0.69fF
C1598 1bitaddie_4/ff_1/m1_58_n52# Gnd 0.24fF
C1599 A4 Gnd 0.55fF
C1600 1bitaddie_4/ff_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1601 1bitaddie_4/ff_0/m1_25_n37# Gnd 0.41fF
C1602 1bitaddie_4/ff_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1603 1bitaddie_4/ff_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1604 1bitaddie_4/ff_0/m1_19_n10# Gnd 0.14fF
C1605 1bitaddie_4/ff_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1606 1bitaddie_4/ff_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1607 1bitaddie_4/ff_0/inverter_0/in Gnd 0.38fF
C1608 1bitaddie_4/ff_0/m1_106_n52# Gnd 0.26fF
C1609 1bitaddie_4/ff_0/m1_63_0# Gnd 0.69fF
C1610 1bitaddie_4/ff_0/m1_58_n52# Gnd 0.24fF
C1611 B4 Gnd 0.61fF
C1612 1bitaddie_4/ff_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1613 1bitaddie_4/xorg_1/m1_102_n17# Gnd 0.04fF
C1614 1bitaddie_4/xorg_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1615 1bitaddie_4/xorg_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1616 1bitaddie_4/xorg_1/m1_25_n11# Gnd 0.13fF
C1617 1bitaddie_4/xorg_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1618 1bitaddie_4/xorg_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1619 1bitaddie_4/xorg_1/m1_102_n91# Gnd 0.22fF
C1620 1bitaddie_4/xorg_1/inverter_1/out Gnd 0.45fF
C1621 1bitaddie_4/sum Gnd 1.47fF
C1622 1bitaddie_4/xorg_1/m1_26_n95# Gnd 0.22fF
C1623 1bitaddie_4/inverter_1/out Gnd 0.90fF
C1624 1bitaddie_4/xorg_1/inverter_1/w_n8_n5# Gnd 0.53fF
C1625 1bitaddie_4/xorg_1/inverter_0/out Gnd 1.68fF
C1626 1bitaddie_4/xorg_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1627 1bitaddie_4/xorg_0/m1_102_n17# Gnd 0.04fF
C1628 1bitaddie_4/xorg_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1629 1bitaddie_4/xorg_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1630 1bitaddie_4/xorg_0/m1_25_n11# Gnd 0.13fF
C1631 1bitaddie_4/xorg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1632 1bitaddie_4/xorg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1633 1bitaddie_4/xorg_0/m1_102_n91# Gnd 0.22fF
C1634 1bitaddie_4/xorg_0/inverter_1/out Gnd 0.45fF
C1635 1bitaddie_4/xorg_0/m1_26_n95# Gnd 0.22fF
C1636 1bitaddie_4/Bi Gnd 1.53fF
C1637 1bitaddie_4/xorg_0/inverter_1/w_n8_n5# Gnd 0.53fF
C1638 1bitaddie_4/xorg_0/inverter_0/out Gnd 1.68fF
C1639 1bitaddie_4/Ai Gnd 2.80fF
C1640 1bitaddie_4/xorg_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1641 inverter_1/out Gnd 3.11fF
C1642 1bitaddie_4/manch_0/clk Gnd 1.66fF
C1643 1bitaddie_4/manch_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1644 1bitaddie_4/manch_0/m1_24_n50# Gnd 0.22fF
C1645 1bitaddie_4/inverter_0/out Gnd 0.59fF
C1646 1bitaddie_4/inverter_2/w_n8_n5# Gnd 0.53fF
C1647 1bitaddie_4/inverter_1/w_n8_n5# Gnd 0.53fF
C1648 1bitaddie_4/inverter_0/w_n8_n5# Gnd 0.53fF
C1649 1bitaddie_4/inverter_0/in Gnd 1.07fF
C1650 1bitaddie_4/nandg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1651 1bitaddie_4/nandg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1652 1bitaddie_4/nandg_0/m1_26_n48# Gnd 0.21fF
C1653 inverter_1/w_n8_n5# Gnd 0.53fF
C1654 inverter_0/in Gnd 0.43fF
C1655 inverter_0/w_n8_n5# Gnd 0.53fF
C1656 1bitaddie_3/Cin Gnd 3.77fF
C1657 1bitaddie_3/ff_2/m1_25_n37# Gnd 0.41fF
C1658 1bitaddie_3/ff_2/pmos_3/w_n8_n5# Gnd 0.58fF
C1659 1bitaddie_3/ff_2/pmos_2/w_n8_n5# Gnd 0.58fF
C1660 1bitaddie_3/ff_2/m1_19_n10# Gnd 0.14fF
C1661 1bitaddie_3/ff_2/pmos_1/w_n8_n5# Gnd 0.58fF
C1662 1bitaddie_3/ff_2/pmos_0/w_n8_n5# Gnd 0.58fF
C1663 1bitaddie_3/ff_2/inverter_0/in Gnd 0.38fF
C1664 1bitaddie_3/ff_2/m1_106_n52# Gnd 0.26fF
C1665 1bitaddie_3/ff_2/m1_63_0# Gnd 0.69fF
C1666 1bitaddie_3/ff_2/m1_58_n52# Gnd 0.24fF
C1667 1bitaddie_3/ff_2/inverter_0/w_n8_n5# Gnd 0.53fF
C1668 1bitaddie_3/ff_1/m1_25_n37# Gnd 0.41fF
C1669 1bitaddie_3/ff_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1670 1bitaddie_3/ff_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1671 1bitaddie_3/ff_1/m1_19_n10# Gnd 0.14fF
C1672 1bitaddie_3/ff_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1673 1bitaddie_3/ff_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1674 1bitaddie_3/ff_1/inverter_0/in Gnd 0.38fF
C1675 1bitaddie_3/ff_1/m1_106_n52# Gnd 0.26fF
C1676 1bitaddie_3/ff_1/m1_63_0# Gnd 0.69fF
C1677 1bitaddie_3/ff_1/m1_58_n52# Gnd 0.24fF
C1678 A3 Gnd 0.55fF
C1679 1bitaddie_3/ff_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1680 1bitaddie_3/ff_0/m1_25_n37# Gnd 0.41fF
C1681 1bitaddie_3/ff_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1682 1bitaddie_3/ff_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1683 1bitaddie_3/ff_0/m1_19_n10# Gnd 0.14fF
C1684 1bitaddie_3/ff_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1685 1bitaddie_3/ff_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1686 1bitaddie_3/ff_0/inverter_0/in Gnd 0.38fF
C1687 1bitaddie_3/ff_0/m1_106_n52# Gnd 0.26fF
C1688 1bitaddie_3/ff_0/m1_63_0# Gnd 0.69fF
C1689 1bitaddie_3/ff_0/m1_58_n52# Gnd 0.24fF
C1690 B3 Gnd 0.61fF
C1691 1bitaddie_3/ff_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1692 1bitaddie_3/xorg_1/m1_102_n17# Gnd 0.04fF
C1693 1bitaddie_3/xorg_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1694 1bitaddie_3/xorg_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1695 1bitaddie_3/xorg_1/m1_25_n11# Gnd 0.13fF
C1696 1bitaddie_3/xorg_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1697 1bitaddie_3/xorg_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1698 1bitaddie_3/xorg_1/m1_102_n91# Gnd 0.22fF
C1699 1bitaddie_3/xorg_1/inverter_1/out Gnd 0.45fF
C1700 1bitaddie_3/sum Gnd 1.47fF
C1701 1bitaddie_3/xorg_1/m1_26_n95# Gnd 0.22fF
C1702 1bitaddie_3/inverter_1/out Gnd 0.90fF
C1703 1bitaddie_3/xorg_1/inverter_1/w_n8_n5# Gnd 0.53fF
C1704 1bitaddie_3/xorg_1/inverter_0/out Gnd 1.68fF
C1705 1bitaddie_3/xorg_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1706 1bitaddie_3/xorg_0/m1_102_n17# Gnd 0.04fF
C1707 1bitaddie_3/xorg_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1708 1bitaddie_3/xorg_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1709 1bitaddie_3/xorg_0/m1_25_n11# Gnd 0.13fF
C1710 1bitaddie_3/xorg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1711 1bitaddie_3/xorg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1712 1bitaddie_3/xorg_0/m1_102_n91# Gnd 0.22fF
C1713 1bitaddie_3/xorg_0/inverter_1/out Gnd 0.45fF
C1714 1bitaddie_3/xorg_0/m1_26_n95# Gnd 0.22fF
C1715 1bitaddie_3/Bi Gnd 1.53fF
C1716 1bitaddie_3/xorg_0/inverter_1/w_n8_n5# Gnd 0.53fF
C1717 1bitaddie_3/xorg_0/inverter_0/out Gnd 1.68fF
C1718 1bitaddie_3/Ai Gnd 2.80fF
C1719 1bitaddie_3/xorg_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1720 1bitaddie_3/manch_0/clk Gnd 1.66fF
C1721 1bitaddie_3/manch_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1722 1bitaddie_3/manch_0/m1_24_n50# Gnd 0.22fF
C1723 1bitaddie_3/inverter_0/out Gnd 0.59fF
C1724 1bitaddie_3/inverter_2/w_n8_n5# Gnd 0.53fF
C1725 1bitaddie_3/inverter_1/w_n8_n5# Gnd 0.53fF
C1726 1bitaddie_3/inverter_0/w_n8_n5# Gnd 0.53fF
C1727 1bitaddie_3/inverter_0/in Gnd 1.07fF
C1728 1bitaddie_3/nandg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1729 1bitaddie_3/nandg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1730 1bitaddie_3/nandg_0/m1_26_n48# Gnd 0.21fF
C1731 1bitaddie_2/Cin Gnd 4.48fF
C1732 1bitaddie_2/ff_2/m1_25_n37# Gnd 0.41fF
C1733 1bitaddie_2/ff_2/pmos_3/w_n8_n5# Gnd 0.58fF
C1734 1bitaddie_2/ff_2/pmos_2/w_n8_n5# Gnd 0.58fF
C1735 1bitaddie_2/ff_2/m1_19_n10# Gnd 0.14fF
C1736 1bitaddie_2/ff_2/pmos_1/w_n8_n5# Gnd 0.58fF
C1737 1bitaddie_2/ff_2/pmos_0/w_n8_n5# Gnd 0.58fF
C1738 1bitaddie_2/ff_2/inverter_0/in Gnd 0.38fF
C1739 1bitaddie_2/ff_2/m1_106_n52# Gnd 0.26fF
C1740 1bitaddie_2/ff_2/m1_63_0# Gnd 0.69fF
C1741 1bitaddie_2/ff_2/m1_58_n52# Gnd 0.24fF
C1742 1bitaddie_2/ff_2/inverter_0/w_n8_n5# Gnd 0.53fF
C1743 1bitaddie_2/ff_1/m1_25_n37# Gnd 0.41fF
C1744 1bitaddie_2/ff_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1745 1bitaddie_2/ff_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1746 1bitaddie_2/ff_1/m1_19_n10# Gnd 0.14fF
C1747 1bitaddie_2/ff_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1748 1bitaddie_2/ff_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1749 1bitaddie_2/ff_1/inverter_0/in Gnd 0.38fF
C1750 1bitaddie_2/ff_1/m1_106_n52# Gnd 0.26fF
C1751 1bitaddie_2/ff_1/m1_63_0# Gnd 0.69fF
C1752 1bitaddie_2/ff_1/m1_58_n52# Gnd 0.24fF
C1753 A2 Gnd 0.55fF
C1754 1bitaddie_2/ff_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1755 1bitaddie_2/ff_0/m1_25_n37# Gnd 0.41fF
C1756 1bitaddie_2/ff_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1757 1bitaddie_2/ff_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1758 1bitaddie_2/ff_0/m1_19_n10# Gnd 0.14fF
C1759 1bitaddie_2/ff_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1760 1bitaddie_2/ff_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1761 1bitaddie_2/ff_0/inverter_0/in Gnd 0.38fF
C1762 1bitaddie_2/ff_0/m1_106_n52# Gnd 0.26fF
C1763 1bitaddie_2/ff_0/m1_63_0# Gnd 0.69fF
C1764 1bitaddie_2/ff_0/m1_58_n52# Gnd 0.24fF
C1765 B2 Gnd 0.61fF
C1766 1bitaddie_2/ff_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1767 1bitaddie_2/xorg_1/m1_102_n17# Gnd 0.04fF
C1768 1bitaddie_2/xorg_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1769 1bitaddie_2/xorg_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1770 1bitaddie_2/xorg_1/m1_25_n11# Gnd 0.13fF
C1771 1bitaddie_2/xorg_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1772 1bitaddie_2/xorg_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1773 1bitaddie_2/xorg_1/m1_102_n91# Gnd 0.22fF
C1774 1bitaddie_2/xorg_1/inverter_1/out Gnd 0.45fF
C1775 1bitaddie_2/sum Gnd 1.47fF
C1776 1bitaddie_2/xorg_1/m1_26_n95# Gnd 0.22fF
C1777 1bitaddie_2/inverter_1/out Gnd 0.90fF
C1778 1bitaddie_2/xorg_1/inverter_1/w_n8_n5# Gnd 0.53fF
C1779 1bitaddie_2/xorg_1/inverter_0/out Gnd 1.68fF
C1780 1bitaddie_2/xorg_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1781 1bitaddie_2/xorg_0/m1_102_n17# Gnd 0.04fF
C1782 1bitaddie_2/xorg_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1783 1bitaddie_2/xorg_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1784 1bitaddie_2/xorg_0/m1_25_n11# Gnd 0.13fF
C1785 1bitaddie_2/xorg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1786 1bitaddie_2/xorg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1787 1bitaddie_2/xorg_0/m1_102_n91# Gnd 0.22fF
C1788 1bitaddie_2/xorg_0/inverter_1/out Gnd 0.45fF
C1789 1bitaddie_2/xorg_0/m1_26_n95# Gnd 0.22fF
C1790 1bitaddie_2/Bi Gnd 1.53fF
C1791 1bitaddie_2/xorg_0/inverter_1/w_n8_n5# Gnd 0.53fF
C1792 1bitaddie_2/xorg_0/inverter_0/out Gnd 1.68fF
C1793 1bitaddie_2/Ai Gnd 2.80fF
C1794 1bitaddie_2/xorg_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1795 1bitaddie_2/manch_0/clk Gnd 1.66fF
C1796 1bitaddie_2/manch_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1797 1bitaddie_2/manch_0/m1_24_n50# Gnd 0.22fF
C1798 1bitaddie_2/inverter_0/out Gnd 0.59fF
C1799 1bitaddie_2/inverter_2/w_n8_n5# Gnd 0.53fF
C1800 1bitaddie_2/inverter_1/w_n8_n5# Gnd 0.53fF
C1801 1bitaddie_2/inverter_0/w_n8_n5# Gnd 0.53fF
C1802 1bitaddie_2/inverter_0/in Gnd 1.07fF
C1803 1bitaddie_2/nandg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1804 1bitaddie_2/nandg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1805 1bitaddie_2/nandg_0/m1_26_n48# Gnd 0.21fF
C1806 1bitaddie_1/Cin Gnd 4.37fF
C1807 1bitaddie_1/ff_2/m1_25_n37# Gnd 0.41fF
C1808 1bitaddie_1/ff_2/pmos_3/w_n8_n5# Gnd 0.58fF
C1809 1bitaddie_1/ff_2/pmos_2/w_n8_n5# Gnd 0.58fF
C1810 1bitaddie_1/ff_2/m1_19_n10# Gnd 0.14fF
C1811 1bitaddie_1/ff_2/pmos_1/w_n8_n5# Gnd 0.58fF
C1812 1bitaddie_1/ff_2/pmos_0/w_n8_n5# Gnd 0.58fF
C1813 1bitaddie_1/ff_2/inverter_0/in Gnd 0.38fF
C1814 1bitaddie_1/ff_2/m1_106_n52# Gnd 0.26fF
C1815 1bitaddie_1/ff_2/m1_63_0# Gnd 0.69fF
C1816 1bitaddie_1/ff_2/m1_58_n52# Gnd 0.24fF
C1817 1bitaddie_1/ff_2/inverter_0/w_n8_n5# Gnd 0.53fF
C1818 1bitaddie_1/ff_1/m1_25_n37# Gnd 0.41fF
C1819 1bitaddie_1/ff_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1820 1bitaddie_1/ff_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1821 1bitaddie_1/ff_1/m1_19_n10# Gnd 0.14fF
C1822 1bitaddie_1/ff_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1823 1bitaddie_1/ff_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1824 1bitaddie_1/ff_1/inverter_0/in Gnd 0.38fF
C1825 1bitaddie_1/ff_1/m1_106_n52# Gnd 0.26fF
C1826 1bitaddie_1/ff_1/m1_63_0# Gnd 0.69fF
C1827 1bitaddie_1/ff_1/m1_58_n52# Gnd 0.24fF
C1828 A1 Gnd 0.55fF
C1829 1bitaddie_1/ff_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1830 1bitaddie_1/ff_0/m1_25_n37# Gnd 0.41fF
C1831 1bitaddie_1/ff_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1832 1bitaddie_1/ff_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1833 1bitaddie_1/ff_0/m1_19_n10# Gnd 0.14fF
C1834 1bitaddie_1/ff_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1835 1bitaddie_1/ff_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1836 1bitaddie_1/ff_0/inverter_0/in Gnd 0.38fF
C1837 1bitaddie_1/ff_0/m1_106_n52# Gnd 0.26fF
C1838 1bitaddie_1/ff_0/m1_63_0# Gnd 0.69fF
C1839 1bitaddie_1/ff_0/m1_58_n52# Gnd 0.24fF
C1840 B1 Gnd 0.60fF
C1841 1bitaddie_1/ff_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1842 1bitaddie_1/xorg_1/m1_102_n17# Gnd 0.04fF
C1843 1bitaddie_1/xorg_1/pmos_3/w_n8_n5# Gnd 0.58fF
C1844 1bitaddie_1/xorg_1/pmos_2/w_n8_n5# Gnd 0.58fF
C1845 1bitaddie_1/xorg_1/m1_25_n11# Gnd 0.13fF
C1846 1bitaddie_1/xorg_1/pmos_1/w_n8_n5# Gnd 0.58fF
C1847 1bitaddie_1/xorg_1/pmos_0/w_n8_n5# Gnd 0.58fF
C1848 1bitaddie_1/xorg_1/m1_102_n91# Gnd 0.22fF
C1849 1bitaddie_1/xorg_1/inverter_1/out Gnd 0.45fF
C1850 1bitaddie_1/sum Gnd 1.47fF
C1851 1bitaddie_1/xorg_1/m1_26_n95# Gnd 0.22fF
C1852 1bitaddie_1/inverter_1/out Gnd 0.90fF
C1853 1bitaddie_1/xorg_1/inverter_1/w_n8_n5# Gnd 0.53fF
C1854 1bitaddie_1/xorg_1/inverter_0/out Gnd 1.68fF
C1855 1bitaddie_1/xorg_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1856 1bitaddie_1/xorg_0/m1_102_n17# Gnd 0.04fF
C1857 1bitaddie_1/xorg_0/pmos_3/w_n8_n5# Gnd 0.58fF
C1858 1bitaddie_1/xorg_0/pmos_2/w_n8_n5# Gnd 0.58fF
C1859 1bitaddie_1/xorg_0/m1_25_n11# Gnd 0.13fF
C1860 1bitaddie_1/xorg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1861 1bitaddie_1/xorg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1862 1bitaddie_1/xorg_0/m1_102_n91# Gnd 0.22fF
C1863 1bitaddie_1/xorg_0/inverter_1/out Gnd 0.45fF
C1864 1bitaddie_1/xorg_0/m1_26_n95# Gnd 0.22fF
C1865 1bitaddie_1/Bi Gnd 1.53fF
C1866 1bitaddie_1/xorg_0/inverter_1/w_n8_n5# Gnd 0.53fF
C1867 1bitaddie_1/xorg_0/inverter_0/out Gnd 1.68fF
C1868 1bitaddie_1/Ai Gnd 2.80fF
C1869 1bitaddie_1/xorg_0/inverter_0/w_n8_n5# Gnd 0.53fF
C1870 1bitaddie_1/manch_0/clk Gnd 1.66fF
C1871 1bitaddie_1/manch_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1872 1bitaddie_1/manch_0/m1_24_n50# Gnd 0.22fF
C1873 1bitaddie_1/inverter_0/out Gnd 0.59fF
C1874 1bitaddie_1/inverter_2/w_n8_n5# Gnd 0.53fF
C1875 1bitaddie_1/inverter_1/w_n8_n5# Gnd 0.53fF
C1876 1bitaddie_1/inverter_0/w_n8_n5# Gnd 0.53fF
C1877 1bitaddie_1/inverter_0/in Gnd 1.07fF
C1878 1bitaddie_1/nandg_0/pmos_1/w_n8_n5# Gnd 0.58fF
C1879 1bitaddie_1/nandg_0/pmos_0/w_n8_n5# Gnd 0.58fF
C1880 1bitaddie_1/nandg_0/m1_26_n48# Gnd 0.21fF

*A0 A1 A2 A3 A4 B0 B1 B2 B3 B4 C0 s0 s1 s2 s3 s4 Cout Vdd Gnd
