magic
tech scmos
timestamp 1764686178
<< nwell >>
rect -5 17 19 40
<< pwell >>
rect -5 -7 19 17
rect -4 -8 19 -7
<< ntransistor >>
rect -34 13 -32 19
rect -18 13 -16 19
rect 6 5 8 11
rect 6 -15 8 -9
<< ptransistor >>
rect 6 23 8 29
<< ndiffusion >>
rect -35 13 -34 19
rect -32 13 -31 19
rect -19 13 -18 19
rect -16 13 -15 19
rect 5 5 6 11
rect 8 5 9 11
rect 5 -15 6 -9
rect 8 -15 9 -9
<< pdiffusion >>
rect 5 23 6 29
rect 8 23 9 29
<< ndcontact >>
rect -39 13 -35 19
rect -31 13 -27 19
rect -23 13 -19 19
rect -15 13 -11 19
rect 1 5 5 11
rect 9 5 13 11
rect 1 -15 5 -9
rect 9 -15 13 -9
<< pdcontact >>
rect 1 23 5 29
rect 9 23 13 29
<< psubstratepcontact >>
rect 9 -3 13 1
rect 1 -23 5 -19
<< nsubstratencontact >>
rect 9 33 13 37
<< polysilicon >>
rect -34 30 8 32
rect -34 19 -32 30
rect 6 29 8 30
rect 6 22 8 23
rect -18 19 -16 22
rect -4 20 8 22
rect -34 6 -32 13
rect -18 6 -16 13
rect -4 -6 -2 20
rect 6 11 8 14
rect 6 -2 8 5
rect -4 -8 8 -6
rect 6 -9 8 -8
rect 6 -18 8 -15
<< polycontact >>
rect -32 6 -28 10
rect -16 6 -12 10
rect 2 -2 6 2
<< metal1 >>
rect 9 29 13 33
rect 1 19 5 23
rect -27 13 -23 19
rect -11 15 25 19
rect -11 13 5 15
rect 1 11 5 13
rect 9 1 13 5
rect 9 -9 13 -3
rect 1 -19 5 -15
<< labels >>
rlabel ndcontact -39 13 -35 19 7 Cc
port 1 w
rlabel polycontact -32 6 -28 10 5 clk
port 2 s
rlabel polycontact -16 6 -12 10 5 P
port 3 s
rlabel polycontact 2 -2 6 2 7 G
port 4 w
rlabel metal1 -11 15 19 19 3 Coc
port 5 e
rlabel psubstratepcontact 1 -23 5 -19 5 gnd
port 6 s
rlabel nsubstratencontact 9 33 13 37 1 vdd
port 7 n
<< end >>
