magic
tech scmos
timestamp 1764797379
<< metal1 >>
rect 118 178 174 183
rect 164 86 172 178
rect 11 77 172 86
rect 53 20 60 41
rect 53 19 100 20
rect 30 15 100 19
rect 44 14 100 15
rect -17 0 3 4
rect 44 -15 50 14
rect 45 -37 50 -15
rect 45 -67 49 -53
rect 45 -97 50 -81
<< m2contact >>
rect 0 77 11 86
rect -6 14 0 19
<< metal2 >>
rect -6 19 0 86
use nmos  nmos_0
timestamp 1764668464
transform 1 0 10 0 1 25
box -10 -25 20 -5
use nmos  nmos_1
timestamp 1764668464
transform 1 0 38 0 1 -30
box -10 -25 20 -5
use nmos  nmos_2
timestamp 1764668464
transform 1 0 38 0 1 -58
box -10 -25 20 -5
use nmos  nmos_3
timestamp 1764668464
transform 1 0 38 0 1 -89
box -10 -25 20 -5
use pmos  pmos_0
timestamp 1764668421
transform 1 0 43 0 1 49
box -10 -11 20 18
use xorg  xorg_0
timestamp 1764782750
transform 1 0 -9 0 1 224
box -62 -125 143 29
<< end >>
