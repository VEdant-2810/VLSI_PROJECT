magic
tech scmos
timestamp 1764813733
<< metal1 >>
rect 648 958 788 961
rect 408 954 488 958
rect 511 955 788 958
rect 408 834 416 954
rect 777 951 788 955
rect 937 953 1164 955
rect 801 950 1164 953
rect 937 946 1164 950
rect 1319 945 1551 946
rect 1184 944 1551 945
rect 1184 942 1555 944
rect 1319 940 1555 942
rect 524 926 527 933
rect 651 927 676 933
rect 815 920 818 925
rect 941 922 957 926
rect 447 907 480 913
rect 572 908 575 915
rect 1197 914 1200 919
rect 1324 915 1339 920
rect 750 900 770 905
rect 862 902 865 907
rect 1245 896 1248 901
rect 486 888 489 895
rect 777 883 780 888
rect 1124 887 1152 893
rect 1159 876 1162 881
rect 522 869 525 876
rect 812 865 815 870
rect 507 858 585 861
rect 589 854 779 859
rect 1195 858 1198 863
rect 796 853 874 856
rect 886 854 1140 857
rect 1137 851 1140 854
rect 1137 847 1165 851
rect 1178 848 1256 851
rect 1271 847 1366 851
rect 67 830 152 834
rect 155 830 417 834
rect 1125 824 1352 825
rect 642 816 715 821
rect 736 816 980 819
rect 1125 817 1362 824
rect 1379 818 1389 940
rect 1536 939 1555 940
rect 1561 936 1698 939
rect 1579 908 1582 913
rect 1703 908 1721 912
rect 1625 890 1628 895
rect 1503 885 1531 890
rect 1541 870 1544 875
rect 1576 852 1579 857
rect 1530 840 1541 843
rect 1556 841 1634 844
rect 642 811 647 816
rect 872 815 980 816
rect 997 815 1362 817
rect 1373 815 1510 818
rect 997 814 1169 815
rect 1133 813 1169 814
rect 80 802 83 807
rect 207 803 218 807
rect 293 801 297 807
rect 420 802 429 806
rect 510 808 647 811
rect 11 780 35 787
rect 127 784 130 792
rect 341 782 345 788
rect 750 787 753 792
rect 877 788 898 792
rect 1012 784 1015 789
rect 1139 786 1153 790
rect 522 779 525 784
rect 649 780 661 784
rect 228 773 248 779
rect 42 762 45 770
rect 255 763 259 769
rect 798 768 801 773
rect 1060 767 1063 772
rect 570 761 573 766
rect 456 756 477 760
rect 672 758 705 765
rect 944 759 968 766
rect 78 744 84 754
rect 292 744 296 750
rect 712 748 715 753
rect 484 742 487 747
rect 974 746 977 751
rect -253 735 44 739
rect 62 735 140 738
rect 150 735 259 738
rect 278 735 356 738
rect -253 725 -244 735
rect 366 734 464 738
rect -253 377 -245 725
rect 461 715 464 734
rect 748 731 751 736
rect 520 724 523 729
rect 1010 728 1013 733
rect 1162 725 1176 734
rect 715 716 722 724
rect 732 720 810 723
rect 824 720 978 724
rect 1144 723 1176 725
rect 969 719 978 720
rect 996 719 1074 722
rect 1085 719 1176 723
rect 1085 718 1145 719
rect 461 711 490 715
rect 507 712 585 715
rect 595 712 727 716
rect 1298 688 1311 815
rect 1388 788 1391 793
rect 1514 788 1526 792
rect 1438 769 1441 774
rect 1316 763 1343 769
rect 1350 749 1353 754
rect 1386 732 1389 737
rect 1637 724 1644 843
rect 1341 707 1351 724
rect 1367 721 1445 724
rect 1460 721 1644 724
rect 1460 720 1634 721
rect 263 619 269 671
rect 550 620 556 676
rect 845 616 854 673
rect 1144 619 1149 672
rect 1463 623 1469 683
rect -32 501 -28 502
rect -32 498 40 501
rect -165 468 -47 471
rect -32 467 -28 498
rect -1 460 8 473
rect 1629 449 1681 453
rect -152 440 -149 445
rect -25 441 -17 445
rect -104 423 -101 428
rect -222 416 -197 422
rect -189 401 -186 406
rect -154 385 -151 390
rect 1674 388 1681 449
rect 1739 436 1955 439
rect 1876 434 1955 436
rect 1756 408 1759 413
rect 1881 409 1917 414
rect 1802 390 1805 395
rect 1674 383 1710 388
rect -253 371 -188 377
rect -168 374 -78 377
rect -97 202 -91 374
rect 1718 369 1721 374
rect 1752 353 1755 358
rect 1735 341 1813 344
rect 1794 328 1802 341
rect 1948 275 1954 434
rect 1750 274 1955 275
rect 1749 269 1955 274
rect 1749 268 1760 269
rect -97 192 21 202
rect -97 -108 -91 192
rect 1554 153 1574 155
rect 1468 150 1574 153
rect 1749 152 1757 268
rect 1554 147 1574 150
rect 1717 148 1766 152
rect 1559 146 1565 147
rect 1580 145 1766 148
rect 1597 117 1600 122
rect 1722 116 1757 121
rect 1645 98 1648 103
rect 278 -57 283 86
rect 340 -16 477 -13
rect 353 -45 356 -40
rect 480 -44 516 -40
rect 278 -64 307 -57
rect 401 -64 404 -59
rect 580 -67 586 82
rect 637 -14 774 -11
rect 653 -42 656 -37
rect 778 -42 803 -37
rect 700 -60 703 -55
rect 916 -67 925 89
rect 959 -4 963 2
rect 983 -7 1120 -4
rect 997 -35 1001 -30
rect 1123 -34 1151 -30
rect 1197 -48 1203 84
rect 1490 79 1550 86
rect 1557 77 1560 82
rect 1596 61 1599 66
rect 1240 -9 1379 -6
rect 1378 -12 1379 -9
rect 1257 -38 1260 -33
rect 1381 -37 1417 -32
rect 1044 -54 1047 -49
rect 1197 -53 1208 -48
rect 1303 -57 1306 -52
rect 580 -74 605 -67
rect 916 -73 951 -67
rect 916 -74 925 -73
rect 960 -74 963 -69
rect 319 -83 322 -78
rect 614 -81 617 -76
rect 1216 -77 1219 -72
rect 995 -92 998 -87
rect 351 -101 354 -96
rect 650 -98 653 -93
rect 1252 -94 1255 -89
rect 636 -108 714 -106
rect 960 -107 965 -100
rect 981 -101 1059 -98
rect 1070 -102 1221 -98
rect 1558 -100 1563 52
rect 1582 50 1660 53
rect 1795 52 1802 230
rect 1669 49 1802 52
rect 1214 -105 1221 -102
rect 1239 -105 1317 -102
rect 1328 -105 1564 -100
rect 722 -108 966 -107
rect -97 -109 317 -108
rect -96 -111 317 -109
rect 339 -112 417 -109
rect 426 -111 966 -108
<< m2contact >>
rect 676 924 686 934
rect 957 918 965 928
rect 1339 912 1350 923
rect 1359 838 1366 847
rect 1721 902 1732 915
rect 1523 838 1530 843
rect 213 798 218 803
rect 429 801 438 810
rect 898 786 906 795
rect 661 777 668 784
rect 1153 782 1160 790
rect 1176 724 1190 734
rect 1526 783 1537 794
rect 1325 707 1341 716
rect 1463 683 1470 688
rect 263 671 269 681
rect 550 676 557 683
rect 845 673 854 681
rect 1144 672 1151 680
rect -24 434 -17 441
rect 1794 318 1800 328
rect 1794 230 1802 241
rect 1766 146 1778 156
rect 477 -21 497 -11
rect 605 -13 614 -1
rect 774 -17 783 -5
rect 945 -5 959 2
rect 1120 -10 1128 -4
rect 1210 -10 1217 -4
rect 1379 -11 1384 -6
<< metal2 >>
rect 213 760 218 798
rect 213 644 217 760
rect 429 711 437 801
rect 263 702 435 711
rect 661 710 666 777
rect 501 707 666 710
rect 263 681 270 702
rect 501 660 505 707
rect 686 703 693 933
rect 957 886 965 918
rect 911 878 965 886
rect 1341 879 1347 912
rect 1302 878 1348 879
rect 911 819 919 878
rect 1297 874 1348 878
rect 1297 873 1322 874
rect 899 718 904 786
rect 550 699 693 703
rect 796 714 904 718
rect 550 683 555 699
rect 796 657 799 714
rect 845 703 851 704
rect 911 703 919 815
rect 1154 760 1158 782
rect 1126 755 1158 760
rect 1126 719 1131 755
rect 1190 725 1204 734
rect 1297 719 1304 873
rect 1366 838 1523 843
rect 1094 718 1131 719
rect 1222 718 1304 719
rect 1091 715 1131 718
rect 845 697 920 703
rect 845 681 851 697
rect 1091 652 1095 715
rect 1126 714 1131 715
rect 1145 715 1304 718
rect 1145 714 1297 715
rect 1145 713 1227 714
rect 1145 680 1152 713
rect 1318 707 1325 717
rect 1464 714 1471 715
rect 1527 714 1533 783
rect 1415 712 1533 714
rect 1412 709 1533 712
rect 1545 776 1551 777
rect 1720 776 1729 902
rect 1545 768 1637 776
rect 1644 768 1730 776
rect 1412 662 1415 709
rect 1545 702 1551 768
rect 1464 699 1551 702
rect 1464 688 1471 699
rect -17 434 -10 441
rect 1794 241 1799 318
rect 497 -17 605 -9
rect 783 -11 952 -5
rect 1128 -9 1210 -5
rect 1766 -7 1777 146
rect 1745 -8 1779 -7
rect 1384 -10 1779 -8
rect 1384 -11 1750 -10
<< m3contact >>
rect 1204 726 1218 734
rect 1318 717 1325 727
rect -10 434 -3 441
<< metal3 >>
rect 1277 734 1331 736
rect 1218 727 1331 734
rect 98 459 101 472
rect -9 445 100 451
rect -9 441 -2 445
use ff  ff_0
timestamp 1764783751
transform 1 0 1721 0 1 412
box -14 -71 160 28
use ff  ff_1
timestamp 1764783751
transform 1 0 1562 0 1 120
box -14 -71 160 28
use ff  ff_2
timestamp 1764783751
transform 1 0 1221 0 1 -34
box -14 -71 160 28
use ff  ff_3
timestamp 1764783751
transform 1 0 963 0 1 -31
box -14 -71 160 28
use ff  ff_4
timestamp 1764783751
transform 1 0 618 0 1 -38
box -14 -71 160 28
use ff  ff_5
timestamp 1764783751
transform 1 0 320 0 1 -41
box -14 -71 160 28
use ff  ff_6
timestamp 1764783751
transform 1 0 -185 0 1 444
box -14 -71 160 28
use ff  ff_7
timestamp 1764783751
transform 1 0 47 0 1 806
box -14 -71 160 28
use ff  ff_8
timestamp 1764783751
transform 1 0 260 0 1 805
box -14 -71 160 28
use ff  ff_10
timestamp 1764783751
transform 1 0 491 0 1 930
box -14 -71 160 28
use ff  ff_9
timestamp 1764783751
transform 1 0 489 0 1 783
box -14 -71 160 28
use ff  ff_12
timestamp 1764783751
transform 1 0 781 0 1 925
box -14 -71 160 28
use ff  ff_11
timestamp 1764783751
transform 1 0 717 0 1 791
box -14 -71 160 28
use ff  ff_13
timestamp 1764783751
transform 1 0 979 0 1 789
box -14 -71 160 28
use ff  ff_14
timestamp 1764783751
transform 1 0 1164 0 1 918
box -14 -71 160 28
use ff  ff_15
timestamp 1764783751
transform 1 0 1354 0 1 791
box -14 -71 160 28
use ff  ff_16
timestamp 1764783751
transform 1 0 1543 0 1 911
box -14 -71 160 28
use cla5_final_without_ff  cla5_final_without_ff_0
timestamp 1764806552
transform 1 0 178 0 1 334
box -178 -334 1472 366
<< labels >>
rlabel metal1 1904 410 1909 411 1 Cout_f
rlabel metal1 1743 116 1750 118 1 S4_f
rlabel metal1 1401 -36 1404 -34 1 S3_f
rlabel metal1 1135 -34 1138 -33 1 S2_f
rlabel metal1 793 -42 797 -40 1 S1_f
rlabel metal1 499 -44 502 -42 1 S0_f
rlabel metal1 -221 416 -218 419 3 Cin_in
rlabel metal1 14 780 17 783 1 A0_in
rlabel metal1 452 907 455 910 1 B1_in
rlabel metal1 459 757 462 758 1 A1_in
rlabel metal1 676 759 681 761 1 A2_in
rlabel metal1 751 901 756 903 1 B2_in
rlabel metal1 947 760 949 761 1 A3_in
rlabel metal1 1128 888 1134 890 1 B3_in
rlabel metal1 1318 765 1322 766 1 A4_in
rlabel metal1 1508 886 1511 888 1 B4_in
rlabel metal1 42 763 43 765 1 clk
rlabel metal1 80 802 83 807 1 clk
rlabel metal1 80 745 81 747 1 clk
rlabel metal1 128 785 129 787 1 clk
rlabel metal1 256 764 257 765 1 clk
rlabel metal1 295 801 296 802 1 clk
rlabel metal1 342 784 343 785 1 clk
rlabel metal1 294 745 295 746 1 clk
rlabel metal1 487 889 488 890 1 clk
rlabel metal1 525 927 526 928 1 clk
rlabel metal1 523 870 524 871 1 clk
rlabel metal1 573 909 574 910 1 clk
rlabel metal1 -188 401 -187 403 1 clk
rlabel metal1 -151 441 -150 443 1 clk
rlabel metal1 -153 385 -152 387 1 clk
rlabel metal1 -103 423 -102 424 1 clk
rlabel metal1 485 743 486 744 1 clk
rlabel metal1 524 780 525 781 1 clk
rlabel metal1 570 762 571 763 1 clk
rlabel metal1 521 725 522 726 1 clk
rlabel metal1 778 884 779 885 1 clk
rlabel metal1 817 921 818 922 1 clk
rlabel metal1 813 866 814 867 1 clk
rlabel metal1 862 905 863 906 1 clk
rlabel metal1 713 750 714 751 1 clk
rlabel metal1 751 788 752 789 1 clk
rlabel metal1 749 732 750 733 1 clk
rlabel metal1 799 769 800 770 1 clk
rlabel metal1 975 748 976 749 1 clk
rlabel metal1 1013 785 1014 786 1 clk
rlabel metal1 1011 730 1012 731 1 clk
rlabel metal1 1061 768 1062 769 1 clk
rlabel metal1 1160 877 1161 878 1 clk
rlabel metal1 1199 915 1200 916 1 clk
rlabel metal1 1196 859 1197 860 1 clk
rlabel metal1 1246 897 1247 898 1 clk
rlabel metal1 1351 750 1352 751 1 clk
rlabel metal1 1389 789 1390 790 1 clk
rlabel metal1 1388 733 1389 734 1 clk
rlabel metal1 1439 770 1440 771 1 clk
rlabel metal1 1542 871 1543 872 1 clk
rlabel metal1 1580 909 1581 910 1 clk
rlabel metal1 1577 853 1578 854 1 clk
rlabel metal1 1627 891 1628 892 1 clk
rlabel metal1 1719 370 1720 371 1 clk
rlabel metal1 1757 409 1758 410 1 clk
rlabel metal1 1752 353 1753 354 1 clk
rlabel metal1 1803 391 1804 392 1 clk
rlabel metal1 1558 79 1559 80 1 clk
rlabel metal1 1598 118 1599 119 1 clk
rlabel metal1 1597 61 1598 62 1 clk
rlabel metal1 1646 99 1647 100 1 clk
rlabel metal1 962 -72 963 -71 1 clk
rlabel metal1 1305 -55 1306 -54 1 clk
rlabel metal1 1254 -92 1255 -91 1 clk
rlabel metal1 1259 -37 1260 -36 1 clk
rlabel metal1 1217 -76 1218 -75 1 clk
rlabel metal1 1044 -53 1045 -52 1 clk
rlabel metal1 996 -90 997 -89 1 clk
rlabel metal1 998 -34 999 -32 1 clk
rlabel metal1 319 -82 320 -81 1 clk
rlabel metal1 354 -44 355 -43 1 clk
rlabel metal1 352 -101 353 -100 1 clk
rlabel metal1 402 -62 403 -61 1 clk
rlabel metal1 615 -79 616 -78 1 clk
rlabel metal1 651 -97 652 -96 1 clk
rlabel metal1 654 -41 655 -40 1 clk
rlabel metal1 701 -59 702 -58 1 clk
rlabel metal1 2 462 6 468 1 clk
rlabel metal3 99 460 100 461 1 clk_mca
<< end >>
